module sprite_rom
	(
		input wire clk,
		input wire [10:0] row,
		input wire [10:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [10:0] row_reg;
	reg [10:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
































































		if(({row_reg, col_reg}>=22'b0000000000000000000000) && ({row_reg, col_reg}<22'b0000100000000001101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100000000001101011) && ({row_reg, col_reg}<22'b0000100000000111101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000100000000111101101) && ({row_reg, col_reg}<22'b0000100000001010010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100000001010010110) && ({row_reg, col_reg}<22'b0000100000010000011000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000100000010000011000) && ({row_reg, col_reg}<22'b0000100000100001100110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100000100001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0000100000100001100111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=22'b0000100000100001101000) && ({row_reg, col_reg}<22'b0000100000100111110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100000100111110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b0000100000100111110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0000100000100111110011) && ({row_reg, col_reg}<22'b0000100000101010010001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100000101010010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b0000100000101010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0000100000101010010011) && ({row_reg, col_reg}<22'b0000100000110000011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100000110000011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==22'b0000100000110000011100)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0000100000110000011101) && ({row_reg, col_reg}<22'b0000100001000001100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100001000001100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==22'b0000100001000001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0000100001000001100101) && ({row_reg, col_reg}<22'b0000100001000111110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100001000111110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0000100001000111110101) && ({row_reg, col_reg}<22'b0000100001001010001110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100001001010001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000100001001010001111) && ({row_reg, col_reg}<22'b0000100001010000011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100001010000011111)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0000100001010000100000) && ({row_reg, col_reg}<22'b0000100001100001100001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100001100001100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000100001100001100010) && ({row_reg, col_reg}<22'b0000100001100111110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100001100111110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0000100001100111110111) && ({row_reg, col_reg}<22'b0000100001101010001100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100001101010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000100001101010001101) && ({row_reg, col_reg}<22'b0000100001110000100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100001110000100001)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0000100001110000100010) && ({row_reg, col_reg}<22'b0000100010000001100000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100010000001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0000100010000001100001) && ({row_reg, col_reg}<22'b0000100010000111111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100010000111111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000100010000111111001) && ({row_reg, col_reg}<22'b0000100010001010001011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100010001010001011) && ({row_reg, col_reg}<22'b0000100010010000100011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000100010010000100011) && ({row_reg, col_reg}<22'b0000100010100001011111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100010100001011111) && ({row_reg, col_reg}<22'b0000100010100111111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100010100111111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0000100010100111111010) && ({row_reg, col_reg}<22'b0000100010101010001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100010101010001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000100010101010001010) && ({row_reg, col_reg}<22'b0000100010110000100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100010110000100100)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0000100010110000100101) && ({row_reg, col_reg}<22'b0000100011000001011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100011000001011110) && ({row_reg, col_reg}<22'b0000100011000111111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100011000111111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0000100011000111111011) && ({row_reg, col_reg}<22'b0000100011001010001000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100011001010001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000100011001010001001) && ({row_reg, col_reg}<22'b0000100011010000100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100011010000100101)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0000100011010000100110) && ({row_reg, col_reg}<22'b0000100011100001011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100011100001011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000100011100001011101) && ({row_reg, col_reg}<22'b0000100011100111111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100011100111111011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0000100011100111111100) && ({row_reg, col_reg}<22'b0000100011101010000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100011101010000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000100011101010001000) && ({row_reg, col_reg}<22'b0000100011110000100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100011110000100110)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0000100011110000100111) && ({row_reg, col_reg}<22'b0000100100000001011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100100000001011100) && ({row_reg, col_reg}<22'b0000100100000111111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100100000111111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0000100100000111111101) && ({row_reg, col_reg}<22'b0000100100001010000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100100001010000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000100100001010000111) && ({row_reg, col_reg}<22'b0000100100010000100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100100010000100111)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0000100100010000101000) && ({row_reg, col_reg}<22'b0000100100100001011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100100100001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0000100100100001011100) && ({row_reg, col_reg}<22'b0000100100100111111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100100100111111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000100100100111111110) && ({row_reg, col_reg}<22'b0000100100101010000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100100101010000110) && ({row_reg, col_reg}<22'b0000100100110000101000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000100100110000101000) && ({row_reg, col_reg}<22'b0000100101000001011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100101000001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000100101000001011011) && ({row_reg, col_reg}<22'b0000100101000111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0000100101000111111110) && ({row_reg, col_reg}<22'b0000100101001010000101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100101001010000101) && ({row_reg, col_reg}<22'b0000100101010000101001)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000100101010000101001) && ({row_reg, col_reg}<22'b0000100101100001011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100101100001011010) && ({row_reg, col_reg}<22'b0000100101100111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100101100111111110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0000100101100111111111) && ({row_reg, col_reg}<22'b0000100101101010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100101101010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000100101101010000101) && ({row_reg, col_reg}<22'b0000100101110000101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100101110000101001)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0000100101110000101010) && ({row_reg, col_reg}<22'b0000100110000001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100110000001011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0000100110000001011010) && ({row_reg, col_reg}<22'b0000100110000111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100110000111111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0000100110001000000000) && ({row_reg, col_reg}<22'b0000100110001010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100110001010000100) && ({row_reg, col_reg}<22'b0000100110010000101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000100110010000101010) && ({row_reg, col_reg}<22'b0000100110100001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100110100001011001) && ({row_reg, col_reg}<22'b0000100110100111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100110100111111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0000100110101000000000) && ({row_reg, col_reg}<22'b0000100110101010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100110101010000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000100110101010000100) && ({row_reg, col_reg}<22'b0000100110110000101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100110110000101010)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0000100110110000101011) && ({row_reg, col_reg}<22'b0000100111000001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000100111000001011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000100111000001011001) && ({row_reg, col_reg}<22'b0000100111001000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100111001000000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000100111001000000001) && ({row_reg, col_reg}<22'b0000100111001010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100111001010000011) && ({row_reg, col_reg}<22'b0000100111010000101011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000100111010000101011) && ({row_reg, col_reg}<22'b0000100111100001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100111100001011000) && ({row_reg, col_reg}<22'b0000100111101000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100111101000000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000100111101000000001) && ({row_reg, col_reg}<22'b0000100111101010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000100111101010000011) && ({row_reg, col_reg}<22'b0000100111110000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000100111110000101011)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000100111110000101100) && ({row_reg, col_reg}<22'b0000101000000001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101000000001011000) && ({row_reg, col_reg}<22'b0000101000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0000101000001000000001) && ({row_reg, col_reg}<22'b0000101000001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101000001010000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101000001010000011) && ({row_reg, col_reg}<22'b0000101000010000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101000010000101011)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0000101000010000101100) && ({row_reg, col_reg}<22'b0000101000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101000100001010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000101000100001011000) && ({row_reg, col_reg}<22'b0000101000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0000101000101000000001) && ({row_reg, col_reg}<22'b0000101000101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101000101010000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0000101000101010000011) && ({row_reg, col_reg}<22'b0000101000110000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101000110000101011)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=22'b0000101000110000101100) && ({row_reg, col_reg}<22'b0000101001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101001000001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0000101001000001011000) && ({row_reg, col_reg}<22'b0000101001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101001001000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101001001000000010) && ({row_reg, col_reg}<22'b0000101001001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101001001010000010) && ({row_reg, col_reg}<22'b0000101001010000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000101001010000101100) && ({row_reg, col_reg}<22'b0000101001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101001100001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0000101001100001011000) && ({row_reg, col_reg}<22'b0000101001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101001101000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000101001101000000010) && ({row_reg, col_reg}<22'b0000101001101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101001101010000010) && ({row_reg, col_reg}<22'b0000101001110000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000101001110000101100) && ({row_reg, col_reg}<22'b0000101010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101010000001010111) && ({row_reg, col_reg}<22'b0000101010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101010001000000010) && ({row_reg, col_reg}<22'b0000101010001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101010001010000010) && ({row_reg, col_reg}<22'b0000101010010000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0000101010010000101100) && ({row_reg, col_reg}<22'b0000101010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101010100001010111) && ({row_reg, col_reg}<22'b0000101010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101010101000000010) && ({row_reg, col_reg}<22'b0000101010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101010101010000010) && ({row_reg, col_reg}<22'b0000101010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101010110000101101) && ({row_reg, col_reg}<22'b0000101011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101011000001010111) && ({row_reg, col_reg}<22'b0000101011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101011001000000010) && ({row_reg, col_reg}<22'b0000101011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101011001010000010) && ({row_reg, col_reg}<22'b0000101011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101011010000101101) && ({row_reg, col_reg}<22'b0000101011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101011100001010111) && ({row_reg, col_reg}<22'b0000101011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101011101000000010) && ({row_reg, col_reg}<22'b0000101011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101011101010000010) && ({row_reg, col_reg}<22'b0000101011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101011110000101101) && ({row_reg, col_reg}<22'b0000101100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101100000001010111) && ({row_reg, col_reg}<22'b0000101100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101100001000000010) && ({row_reg, col_reg}<22'b0000101100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101100001010000010) && ({row_reg, col_reg}<22'b0000101100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101100010000101101) && ({row_reg, col_reg}<22'b0000101100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101100100001010111) && ({row_reg, col_reg}<22'b0000101100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101100101000000010) && ({row_reg, col_reg}<22'b0000101100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101100101010000010) && ({row_reg, col_reg}<22'b0000101100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101100110000101101) && ({row_reg, col_reg}<22'b0000101101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101101000001010111) && ({row_reg, col_reg}<22'b0000101101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101101001000000010) && ({row_reg, col_reg}<22'b0000101101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101101001010000010) && ({row_reg, col_reg}<22'b0000101101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101101010000101101) && ({row_reg, col_reg}<22'b0000101101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101101100001010111) && ({row_reg, col_reg}<22'b0000101101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000101101101000000010) && ({row_reg, col_reg}<22'b0000101101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101101101010000010) && ({row_reg, col_reg}<22'b0000101101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101101110000101101) && ({row_reg, col_reg}<22'b0000101110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101110000001010111) && ({row_reg, col_reg}<22'b0000101110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101110001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000101110001000000010) && ({row_reg, col_reg}<22'b0000101110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101110001010000010) && ({row_reg, col_reg}<22'b0000101110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101110010000101101) && ({row_reg, col_reg}<22'b0000101110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101110100001010111) && ({row_reg, col_reg}<22'b0000101110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000101110101000000010) && ({row_reg, col_reg}<22'b0000101110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101110101010000010) && ({row_reg, col_reg}<22'b0000101110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101110110000101101) && ({row_reg, col_reg}<22'b0000101111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101111000001010111) && ({row_reg, col_reg}<22'b0000101111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101111001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000101111001000000010) && ({row_reg, col_reg}<22'b0000101111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101111001010000010) && ({row_reg, col_reg}<22'b0000101111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101111010000101101) && ({row_reg, col_reg}<22'b0000101111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000101111100001010111) && ({row_reg, col_reg}<22'b0000101111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101111101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000101111101000000010) && ({row_reg, col_reg}<22'b0000101111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000101111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000101111101010000010) && ({row_reg, col_reg}<22'b0000101111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000101111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000101111110000101101) && ({row_reg, col_reg}<22'b0000110000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110000000001010111) && ({row_reg, col_reg}<22'b0000110000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110000001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000110000001000000010) && ({row_reg, col_reg}<22'b0000110000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110000001010000010) && ({row_reg, col_reg}<22'b0000110000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110000010000101101) && ({row_reg, col_reg}<22'b0000110000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110000100001010111) && ({row_reg, col_reg}<22'b0000110000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000110000101000000010) && ({row_reg, col_reg}<22'b0000110000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110000101010000010) && ({row_reg, col_reg}<22'b0000110000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110000110000101101) && ({row_reg, col_reg}<22'b0000110001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110001000001010111) && ({row_reg, col_reg}<22'b0000110001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110001001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000110001001000000010) && ({row_reg, col_reg}<22'b0000110001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110001001010000010) && ({row_reg, col_reg}<22'b0000110001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110001010000101101) && ({row_reg, col_reg}<22'b0000110001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110001100001010111) && ({row_reg, col_reg}<22'b0000110001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110001101000000010) && ({row_reg, col_reg}<22'b0000110001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110001101010000010) && ({row_reg, col_reg}<22'b0000110001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110001110000101101) && ({row_reg, col_reg}<22'b0000110010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110010000001010111) && ({row_reg, col_reg}<22'b0000110010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110010001000000010) && ({row_reg, col_reg}<22'b0000110010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110010001010000010) && ({row_reg, col_reg}<22'b0000110010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110010010000101101) && ({row_reg, col_reg}<22'b0000110010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110010100001010111) && ({row_reg, col_reg}<22'b0000110010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110010101000000010) && ({row_reg, col_reg}<22'b0000110010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110010101010000010) && ({row_reg, col_reg}<22'b0000110010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110010110000101101) && ({row_reg, col_reg}<22'b0000110011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110011000001010111) && ({row_reg, col_reg}<22'b0000110011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110011001000000010) && ({row_reg, col_reg}<22'b0000110011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110011001010000010) && ({row_reg, col_reg}<22'b0000110011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110011010000101101) && ({row_reg, col_reg}<22'b0000110011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110011100001010111) && ({row_reg, col_reg}<22'b0000110011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110011101000000010) && ({row_reg, col_reg}<22'b0000110011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110011101010000010) && ({row_reg, col_reg}<22'b0000110011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110011110000101101) && ({row_reg, col_reg}<22'b0000110100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110100000001010111) && ({row_reg, col_reg}<22'b0000110100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110100001000000010) && ({row_reg, col_reg}<22'b0000110100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110100001010000010) && ({row_reg, col_reg}<22'b0000110100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110100010000101101) && ({row_reg, col_reg}<22'b0000110100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110100100001010111) && ({row_reg, col_reg}<22'b0000110100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110100101000000010) && ({row_reg, col_reg}<22'b0000110100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110100101010000010) && ({row_reg, col_reg}<22'b0000110100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110100110000101101) && ({row_reg, col_reg}<22'b0000110101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110101000001010111) && ({row_reg, col_reg}<22'b0000110101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110101001000000010) && ({row_reg, col_reg}<22'b0000110101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110101001010000010) && ({row_reg, col_reg}<22'b0000110101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110101010000101101) && ({row_reg, col_reg}<22'b0000110101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110101100001010111) && ({row_reg, col_reg}<22'b0000110101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110101100010000001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=22'b0000110101100010000010) && ({row_reg, col_reg}<22'b0000110101100111010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110101100111010111) && ({row_reg, col_reg}<22'b0000110101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110101101000000010) && ({row_reg, col_reg}<22'b0000110101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110101101010000010) && ({row_reg, col_reg}<22'b0000110101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110101101010101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000110101101010101101) && ({row_reg, col_reg}<22'b0000110101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==22'b0000110101110000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0000110101110000000010) && ({row_reg, col_reg}<22'b0000110101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110101110000101101) && ({row_reg, col_reg}<22'b0000110110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110110000001010111) && ({row_reg, col_reg}<22'b0000110110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110110000010000010) && ({row_reg, col_reg}<22'b0000110110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110110000111010111) && ({row_reg, col_reg}<22'b0000110110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110110001000000010) && ({row_reg, col_reg}<22'b0000110110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110110001010000010) && ({row_reg, col_reg}<22'b0000110110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110110001010101101) && ({row_reg, col_reg}<22'b0000110110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110110010000000010) && ({row_reg, col_reg}<22'b0000110110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110110010000101101) && ({row_reg, col_reg}<22'b0000110110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110110100001010111) && ({row_reg, col_reg}<22'b0000110110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110110100010000010) && ({row_reg, col_reg}<22'b0000110110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110110100111010111) && ({row_reg, col_reg}<22'b0000110110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110110101000000010) && ({row_reg, col_reg}<22'b0000110110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110110101010000010) && ({row_reg, col_reg}<22'b0000110110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110110101010101101) && ({row_reg, col_reg}<22'b0000110110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110110110000000010) && ({row_reg, col_reg}<22'b0000110110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110110110000101101) && ({row_reg, col_reg}<22'b0000110111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110111000001010111) && ({row_reg, col_reg}<22'b0000110111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110111000010000010) && ({row_reg, col_reg}<22'b0000110111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110111000111010111) && ({row_reg, col_reg}<22'b0000110111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110111001000000010) && ({row_reg, col_reg}<22'b0000110111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110111001010000010) && ({row_reg, col_reg}<22'b0000110111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110111001010101101) && ({row_reg, col_reg}<22'b0000110111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110111010000000010) && ({row_reg, col_reg}<22'b0000110111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110111010000101101) && ({row_reg, col_reg}<22'b0000110111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110111100001010111) && ({row_reg, col_reg}<22'b0000110111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110111100010000010) && ({row_reg, col_reg}<22'b0000110111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000110111100111010111) && ({row_reg, col_reg}<22'b0000110111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000110111101000000010) && ({row_reg, col_reg}<22'b0000110111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110111101010000010) && ({row_reg, col_reg}<22'b0000110111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110111101010101101) && ({row_reg, col_reg}<22'b0000110111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000110111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000110111110000000010) && ({row_reg, col_reg}<22'b0000110111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000110111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000110111110000101101) && ({row_reg, col_reg}<22'b0000111000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111000000001010111) && ({row_reg, col_reg}<22'b0000111000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111000000010000010) && ({row_reg, col_reg}<22'b0000111000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111000000111010111) && ({row_reg, col_reg}<22'b0000111000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111000001000000010) && ({row_reg, col_reg}<22'b0000111000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111000001010000010) && ({row_reg, col_reg}<22'b0000111000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111000001010101101) && ({row_reg, col_reg}<22'b0000111000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111000010000000010) && ({row_reg, col_reg}<22'b0000111000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111000010000101101) && ({row_reg, col_reg}<22'b0000111000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111000100001010111) && ({row_reg, col_reg}<22'b0000111000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111000100010000010) && ({row_reg, col_reg}<22'b0000111000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111000100111010111) && ({row_reg, col_reg}<22'b0000111000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111000101000000010) && ({row_reg, col_reg}<22'b0000111000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111000101010000010) && ({row_reg, col_reg}<22'b0000111000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111000101010101101) && ({row_reg, col_reg}<22'b0000111000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111000110000000010) && ({row_reg, col_reg}<22'b0000111000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111000110000101101) && ({row_reg, col_reg}<22'b0000111001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111001000001010111) && ({row_reg, col_reg}<22'b0000111001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111001000010000010) && ({row_reg, col_reg}<22'b0000111001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111001000111010111) && ({row_reg, col_reg}<22'b0000111001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000111001001000000010) && ({row_reg, col_reg}<22'b0000111001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111001001010000010) && ({row_reg, col_reg}<22'b0000111001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111001001010101101) && ({row_reg, col_reg}<22'b0000111001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111001010000000010) && ({row_reg, col_reg}<22'b0000111001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111001010000101101) && ({row_reg, col_reg}<22'b0000111001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111001100001010111) && ({row_reg, col_reg}<22'b0000111001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111001100010000010) && ({row_reg, col_reg}<22'b0000111001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111001100111010111) && ({row_reg, col_reg}<22'b0000111001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000111001101000000010) && ({row_reg, col_reg}<22'b0000111001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111001101010000010) && ({row_reg, col_reg}<22'b0000111001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111001101010101101) && ({row_reg, col_reg}<22'b0000111001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111001110000000010) && ({row_reg, col_reg}<22'b0000111001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111001110000101101) && ({row_reg, col_reg}<22'b0000111010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111010000001010111) && ({row_reg, col_reg}<22'b0000111010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111010000010000010) && ({row_reg, col_reg}<22'b0000111010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111010000111010111) && ({row_reg, col_reg}<22'b0000111010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000111010001000000010) && ({row_reg, col_reg}<22'b0000111010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111010001010000010) && ({row_reg, col_reg}<22'b0000111010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111010001010101101) && ({row_reg, col_reg}<22'b0000111010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111010010000000010) && ({row_reg, col_reg}<22'b0000111010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111010010000101101) && ({row_reg, col_reg}<22'b0000111010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111010100001010111) && ({row_reg, col_reg}<22'b0000111010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111010100010000010) && ({row_reg, col_reg}<22'b0000111010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111010100111010111) && ({row_reg, col_reg}<22'b0000111010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111010101000000010) && ({row_reg, col_reg}<22'b0000111010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111010101010000010) && ({row_reg, col_reg}<22'b0000111010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111010101010101101) && ({row_reg, col_reg}<22'b0000111010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111010110000000010) && ({row_reg, col_reg}<22'b0000111010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111010110000101101) && ({row_reg, col_reg}<22'b0000111011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111011000001010111) && ({row_reg, col_reg}<22'b0000111011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000111011000010000010) && ({row_reg, col_reg}<22'b0000111011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111011000111010111) && ({row_reg, col_reg}<22'b0000111011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111011001000000010) && ({row_reg, col_reg}<22'b0000111011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111011001010000010) && ({row_reg, col_reg}<22'b0000111011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111011001010101101) && ({row_reg, col_reg}<22'b0000111011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111011010000000010) && ({row_reg, col_reg}<22'b0000111011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111011010000101101) && ({row_reg, col_reg}<22'b0000111011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111011100001010111) && ({row_reg, col_reg}<22'b0000111011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000111011100010000010) && ({row_reg, col_reg}<22'b0000111011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111011100111010111) && ({row_reg, col_reg}<22'b0000111011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111011101000000010) && ({row_reg, col_reg}<22'b0000111011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111011101010000010) && ({row_reg, col_reg}<22'b0000111011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111011101010101101) && ({row_reg, col_reg}<22'b0000111011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111011110000000010) && ({row_reg, col_reg}<22'b0000111011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111011110000101101) && ({row_reg, col_reg}<22'b0000111100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111100000001010111) && ({row_reg, col_reg}<22'b0000111100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0000111100000010000010) && ({row_reg, col_reg}<22'b0000111100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111100000111010111) && ({row_reg, col_reg}<22'b0000111100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111100001000000010) && ({row_reg, col_reg}<22'b0000111100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111100001010000010) && ({row_reg, col_reg}<22'b0000111100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111100001010101101) && ({row_reg, col_reg}<22'b0000111100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111100010000000010) && ({row_reg, col_reg}<22'b0000111100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111100010000101101) && ({row_reg, col_reg}<22'b0000111100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111100100001010111) && ({row_reg, col_reg}<22'b0000111100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111100100010000010) && ({row_reg, col_reg}<22'b0000111100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111100100111010111) && ({row_reg, col_reg}<22'b0000111100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111100101000000010) && ({row_reg, col_reg}<22'b0000111100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111100101010000010) && ({row_reg, col_reg}<22'b0000111100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111100101010101101) && ({row_reg, col_reg}<22'b0000111100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111100110000000010) && ({row_reg, col_reg}<22'b0000111100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111100110000101101) && ({row_reg, col_reg}<22'b0000111101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111101000001010111) && ({row_reg, col_reg}<22'b0000111101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0000111101000010000010) && ({row_reg, col_reg}<22'b0000111101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111101000111010111) && ({row_reg, col_reg}<22'b0000111101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111101001000000010) && ({row_reg, col_reg}<22'b0000111101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111101001010000010) && ({row_reg, col_reg}<22'b0000111101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111101001010101101) && ({row_reg, col_reg}<22'b0000111101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111101010000000010) && ({row_reg, col_reg}<22'b0000111101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111101010000101101) && ({row_reg, col_reg}<22'b0000111101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111101100001010111) && ({row_reg, col_reg}<22'b0000111101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111101100010000010) && ({row_reg, col_reg}<22'b0000111101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111101100111010111) && ({row_reg, col_reg}<22'b0000111101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111101101000000010) && ({row_reg, col_reg}<22'b0000111101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111101101010000010) && ({row_reg, col_reg}<22'b0000111101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111101101010101101) && ({row_reg, col_reg}<22'b0000111101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111101110000000010) && ({row_reg, col_reg}<22'b0000111101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111101110000101101) && ({row_reg, col_reg}<22'b0000111110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111110000001010111) && ({row_reg, col_reg}<22'b0000111110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111110000010000010) && ({row_reg, col_reg}<22'b0000111110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111110000111010111) && ({row_reg, col_reg}<22'b0000111110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111110001000000010) && ({row_reg, col_reg}<22'b0000111110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111110001010000010) && ({row_reg, col_reg}<22'b0000111110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111110001010101101) && ({row_reg, col_reg}<22'b0000111110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111110010000000010) && ({row_reg, col_reg}<22'b0000111110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111110010000101101) && ({row_reg, col_reg}<22'b0000111110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111110100001010111) && ({row_reg, col_reg}<22'b0000111110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111110100010000010) && ({row_reg, col_reg}<22'b0000111110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111110100111010111) && ({row_reg, col_reg}<22'b0000111110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111110101000000010) && ({row_reg, col_reg}<22'b0000111110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111110101010000010) && ({row_reg, col_reg}<22'b0000111110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111110101010101101) && ({row_reg, col_reg}<22'b0000111110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111110110000000010) && ({row_reg, col_reg}<22'b0000111110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111110110000101101) && ({row_reg, col_reg}<22'b0000111111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111111000001010111) && ({row_reg, col_reg}<22'b0000111111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111111000010000010) && ({row_reg, col_reg}<22'b0000111111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111111000111010111) && ({row_reg, col_reg}<22'b0000111111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111111001000000010) && ({row_reg, col_reg}<22'b0000111111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111111001010000010) && ({row_reg, col_reg}<22'b0000111111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111111001010101101) && ({row_reg, col_reg}<22'b0000111111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111111010000000010) && ({row_reg, col_reg}<22'b0000111111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111111010000101101) && ({row_reg, col_reg}<22'b0000111111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111111100001010111) && ({row_reg, col_reg}<22'b0000111111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111111100010000010) && ({row_reg, col_reg}<22'b0000111111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0000111111100111010111) && ({row_reg, col_reg}<22'b0000111111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0000111111101000000010) && ({row_reg, col_reg}<22'b0000111111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111111101010000010) && ({row_reg, col_reg}<22'b0000111111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111111101010101101) && ({row_reg, col_reg}<22'b0000111111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0000111111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0000111111110000000010) && ({row_reg, col_reg}<22'b0000111111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0000111111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0000111111110000101101) && ({row_reg, col_reg}<22'b0001000000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000000000001010111) && ({row_reg, col_reg}<22'b0001000000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000000000010000010) && ({row_reg, col_reg}<22'b0001000000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000000000111010111) && ({row_reg, col_reg}<22'b0001000000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000000001000000010) && ({row_reg, col_reg}<22'b0001000000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000000001010000010) && ({row_reg, col_reg}<22'b0001000000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000000001010101101) && ({row_reg, col_reg}<22'b0001000000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000000010000000010) && ({row_reg, col_reg}<22'b0001000000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000000010000101101) && ({row_reg, col_reg}<22'b0001000000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000000100001010111) && ({row_reg, col_reg}<22'b0001000000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000000100010000010) && ({row_reg, col_reg}<22'b0001000000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000000100111010111) && ({row_reg, col_reg}<22'b0001000000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000000101000000010) && ({row_reg, col_reg}<22'b0001000000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000000101010000010) && ({row_reg, col_reg}<22'b0001000000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000000101010101101) && ({row_reg, col_reg}<22'b0001000000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000000110000000010) && ({row_reg, col_reg}<22'b0001000000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000000110000101101) && ({row_reg, col_reg}<22'b0001000001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000001000001010111) && ({row_reg, col_reg}<22'b0001000001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000001000010000010) && ({row_reg, col_reg}<22'b0001000001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000001000111010111) && ({row_reg, col_reg}<22'b0001000001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000001001000000010) && ({row_reg, col_reg}<22'b0001000001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000001001010000010) && ({row_reg, col_reg}<22'b0001000001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000001001010101101) && ({row_reg, col_reg}<22'b0001000001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000001010000000010) && ({row_reg, col_reg}<22'b0001000001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000001010000101101) && ({row_reg, col_reg}<22'b0001000001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000001100001010111) && ({row_reg, col_reg}<22'b0001000001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000001100010000010) && ({row_reg, col_reg}<22'b0001000001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000001100111010111) && ({row_reg, col_reg}<22'b0001000001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000001101000000010) && ({row_reg, col_reg}<22'b0001000001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000001101010000010) && ({row_reg, col_reg}<22'b0001000001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000001101010101101) && ({row_reg, col_reg}<22'b0001000001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000001110000000010) && ({row_reg, col_reg}<22'b0001000001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000001110000101101) && ({row_reg, col_reg}<22'b0001000010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000010000001010111) && ({row_reg, col_reg}<22'b0001000010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000010000010000010) && ({row_reg, col_reg}<22'b0001000010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000010000111010111) && ({row_reg, col_reg}<22'b0001000010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000010001000000010) && ({row_reg, col_reg}<22'b0001000010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000010001010000010) && ({row_reg, col_reg}<22'b0001000010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000010001010101101) && ({row_reg, col_reg}<22'b0001000010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000010010000000010) && ({row_reg, col_reg}<22'b0001000010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000010010000101101) && ({row_reg, col_reg}<22'b0001000010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000010100001010111) && ({row_reg, col_reg}<22'b0001000010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000010100010000010) && ({row_reg, col_reg}<22'b0001000010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000010100111010111) && ({row_reg, col_reg}<22'b0001000010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000010101000000010) && ({row_reg, col_reg}<22'b0001000010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000010101010000010) && ({row_reg, col_reg}<22'b0001000010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000010101010101101) && ({row_reg, col_reg}<22'b0001000010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000010110000000010) && ({row_reg, col_reg}<22'b0001000010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000010110000101101) && ({row_reg, col_reg}<22'b0001000011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000011000001010111) && ({row_reg, col_reg}<22'b0001000011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000011000010000010) && ({row_reg, col_reg}<22'b0001000011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000011000111010111) && ({row_reg, col_reg}<22'b0001000011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001000011001000000010) && ({row_reg, col_reg}<22'b0001000011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000011001010000010) && ({row_reg, col_reg}<22'b0001000011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000011001010101101) && ({row_reg, col_reg}<22'b0001000011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000011010000000010) && ({row_reg, col_reg}<22'b0001000011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000011010000101101) && ({row_reg, col_reg}<22'b0001000011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000011100001010111) && ({row_reg, col_reg}<22'b0001000011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000011100010000010) && ({row_reg, col_reg}<22'b0001000011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000011100111010111) && ({row_reg, col_reg}<22'b0001000011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001000011101000000010) && ({row_reg, col_reg}<22'b0001000011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000011101010000010) && ({row_reg, col_reg}<22'b0001000011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000011101010101101) && ({row_reg, col_reg}<22'b0001000011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000011110000000010) && ({row_reg, col_reg}<22'b0001000011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000011110000101101) && ({row_reg, col_reg}<22'b0001000100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000100000001010111) && ({row_reg, col_reg}<22'b0001000100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000100000010000010) && ({row_reg, col_reg}<22'b0001000100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000100000111010111) && ({row_reg, col_reg}<22'b0001000100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001000100001000000010) && ({row_reg, col_reg}<22'b0001000100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000100001010000010) && ({row_reg, col_reg}<22'b0001000100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000100001010101101) && ({row_reg, col_reg}<22'b0001000100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000100010000000010) && ({row_reg, col_reg}<22'b0001000100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000100010000101101) && ({row_reg, col_reg}<22'b0001000100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000100100001010111) && ({row_reg, col_reg}<22'b0001000100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000100100010000010) && ({row_reg, col_reg}<22'b0001000100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000100100111010111) && ({row_reg, col_reg}<22'b0001000100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000100101000000010) && ({row_reg, col_reg}<22'b0001000100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000100101010000010) && ({row_reg, col_reg}<22'b0001000100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000100101010101101) && ({row_reg, col_reg}<22'b0001000100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000100110000000010) && ({row_reg, col_reg}<22'b0001000100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000100110000101101) && ({row_reg, col_reg}<22'b0001000101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000101000001010111) && ({row_reg, col_reg}<22'b0001000101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001000101000010000010) && ({row_reg, col_reg}<22'b0001000101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000101000111010111) && ({row_reg, col_reg}<22'b0001000101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000101001000000010) && ({row_reg, col_reg}<22'b0001000101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000101001010000010) && ({row_reg, col_reg}<22'b0001000101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000101001010101101) && ({row_reg, col_reg}<22'b0001000101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000101010000000010) && ({row_reg, col_reg}<22'b0001000101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000101010000101101) && ({row_reg, col_reg}<22'b0001000101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000101100001010111) && ({row_reg, col_reg}<22'b0001000101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001000101100010000010) && ({row_reg, col_reg}<22'b0001000101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000101100111010111) && ({row_reg, col_reg}<22'b0001000101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000101101000000010) && ({row_reg, col_reg}<22'b0001000101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000101101010000010) && ({row_reg, col_reg}<22'b0001000101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000101101010101101) && ({row_reg, col_reg}<22'b0001000101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000101110000000010) && ({row_reg, col_reg}<22'b0001000101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000101110000101101) && ({row_reg, col_reg}<22'b0001000110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000110000001010111) && ({row_reg, col_reg}<22'b0001000110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001000110000010000010) && ({row_reg, col_reg}<22'b0001000110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000110000111010111) && ({row_reg, col_reg}<22'b0001000110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000110001000000010) && ({row_reg, col_reg}<22'b0001000110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000110001010000010) && ({row_reg, col_reg}<22'b0001000110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000110001010101101) && ({row_reg, col_reg}<22'b0001000110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000110010000000010) && ({row_reg, col_reg}<22'b0001000110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000110010000101101) && ({row_reg, col_reg}<22'b0001000110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000110100001010111) && ({row_reg, col_reg}<22'b0001000110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000110100010000010) && ({row_reg, col_reg}<22'b0001000110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000110100111010111) && ({row_reg, col_reg}<22'b0001000110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000110101000000010) && ({row_reg, col_reg}<22'b0001000110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000110101010000010) && ({row_reg, col_reg}<22'b0001000110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000110101010101101) && ({row_reg, col_reg}<22'b0001000110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000110110000000010) && ({row_reg, col_reg}<22'b0001000110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000110110000101101) && ({row_reg, col_reg}<22'b0001000111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000111000001010111) && ({row_reg, col_reg}<22'b0001000111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001000111000010000010) && ({row_reg, col_reg}<22'b0001000111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000111000111010111) && ({row_reg, col_reg}<22'b0001000111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000111001000000010) && ({row_reg, col_reg}<22'b0001000111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000111001010000010) && ({row_reg, col_reg}<22'b0001000111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000111001010101101) && ({row_reg, col_reg}<22'b0001000111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000111010000000010) && ({row_reg, col_reg}<22'b0001000111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000111010000101101) && ({row_reg, col_reg}<22'b0001000111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000111100001010111) && ({row_reg, col_reg}<22'b0001000111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000111100010000010) && ({row_reg, col_reg}<22'b0001000111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001000111100111010111) && ({row_reg, col_reg}<22'b0001000111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001000111101000000010) && ({row_reg, col_reg}<22'b0001000111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000111101010000010) && ({row_reg, col_reg}<22'b0001000111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000111101010101101) && ({row_reg, col_reg}<22'b0001000111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001000111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001000111110000000010) && ({row_reg, col_reg}<22'b0001000111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001000111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001000111110000101101) && ({row_reg, col_reg}<22'b0001001000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001000000001010111) && ({row_reg, col_reg}<22'b0001001000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001000000010000010) && ({row_reg, col_reg}<22'b0001001000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001000000111010111) && ({row_reg, col_reg}<22'b0001001000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001000001000000010) && ({row_reg, col_reg}<22'b0001001000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001000001010000010) && ({row_reg, col_reg}<22'b0001001000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001000001010101101) && ({row_reg, col_reg}<22'b0001001000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001000010000000010) && ({row_reg, col_reg}<22'b0001001000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001000010000101101) && ({row_reg, col_reg}<22'b0001001000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001000100001010111) && ({row_reg, col_reg}<22'b0001001000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001000100010000010) && ({row_reg, col_reg}<22'b0001001000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001000100111010111) && ({row_reg, col_reg}<22'b0001001000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001000101000000010) && ({row_reg, col_reg}<22'b0001001000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001000101010000010) && ({row_reg, col_reg}<22'b0001001000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001000101010101101) && ({row_reg, col_reg}<22'b0001001000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001000110000000010) && ({row_reg, col_reg}<22'b0001001000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001000110000101101) && ({row_reg, col_reg}<22'b0001001001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001001000001010111) && ({row_reg, col_reg}<22'b0001001001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001001000010000010) && ({row_reg, col_reg}<22'b0001001001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001001000111010111) && ({row_reg, col_reg}<22'b0001001001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001001001000000010) && ({row_reg, col_reg}<22'b0001001001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001001001010000010) && ({row_reg, col_reg}<22'b0001001001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001001001010101101) && ({row_reg, col_reg}<22'b0001001001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001001010000000010) && ({row_reg, col_reg}<22'b0001001001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001001010000101101) && ({row_reg, col_reg}<22'b0001001001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001001100001010111) && ({row_reg, col_reg}<22'b0001001001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001001100010000010) && ({row_reg, col_reg}<22'b0001001001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001001100111010111) && ({row_reg, col_reg}<22'b0001001001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001001101000000010) && ({row_reg, col_reg}<22'b0001001001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001001101010000010) && ({row_reg, col_reg}<22'b0001001001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001001101010101101) && ({row_reg, col_reg}<22'b0001001001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001001110000000010) && ({row_reg, col_reg}<22'b0001001001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001001110000101101) && ({row_reg, col_reg}<22'b0001001010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001010000001010111) && ({row_reg, col_reg}<22'b0001001010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001010000010000010) && ({row_reg, col_reg}<22'b0001001010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001010000111010111) && ({row_reg, col_reg}<22'b0001001010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001010001000000010) && ({row_reg, col_reg}<22'b0001001010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001010001010000010) && ({row_reg, col_reg}<22'b0001001010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001010001010101101) && ({row_reg, col_reg}<22'b0001001010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001010010000000010) && ({row_reg, col_reg}<22'b0001001010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001010010000101101) && ({row_reg, col_reg}<22'b0001001010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001010100001010111) && ({row_reg, col_reg}<22'b0001001010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001010100010000010) && ({row_reg, col_reg}<22'b0001001010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001010100111010111) && ({row_reg, col_reg}<22'b0001001010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001010101000000010) && ({row_reg, col_reg}<22'b0001001010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001010101010000010) && ({row_reg, col_reg}<22'b0001001010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001010101010101101) && ({row_reg, col_reg}<22'b0001001010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001010110000000010) && ({row_reg, col_reg}<22'b0001001010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001010110000101101) && ({row_reg, col_reg}<22'b0001001011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001011000001010111) && ({row_reg, col_reg}<22'b0001001011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001011000010000010) && ({row_reg, col_reg}<22'b0001001011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001011000111010111) && ({row_reg, col_reg}<22'b0001001011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001011001000000010) && ({row_reg, col_reg}<22'b0001001011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001011001010000010) && ({row_reg, col_reg}<22'b0001001011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001011001010101101) && ({row_reg, col_reg}<22'b0001001011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001011010000000010) && ({row_reg, col_reg}<22'b0001001011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001011010000101101) && ({row_reg, col_reg}<22'b0001001011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001011100001010111) && ({row_reg, col_reg}<22'b0001001011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001011100010000010) && ({row_reg, col_reg}<22'b0001001011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001011100111010111) && ({row_reg, col_reg}<22'b0001001011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001011101000000010) && ({row_reg, col_reg}<22'b0001001011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001011101010000010) && ({row_reg, col_reg}<22'b0001001011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001011101010101101) && ({row_reg, col_reg}<22'b0001001011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001011110000000010) && ({row_reg, col_reg}<22'b0001001011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001011110000101101) && ({row_reg, col_reg}<22'b0001001100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001100000001010111) && ({row_reg, col_reg}<22'b0001001100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001100000010000010) && ({row_reg, col_reg}<22'b0001001100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001100000111010111) && ({row_reg, col_reg}<22'b0001001100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001001100001000000010) && ({row_reg, col_reg}<22'b0001001100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001100001010000010) && ({row_reg, col_reg}<22'b0001001100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001100001010101101) && ({row_reg, col_reg}<22'b0001001100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001100010000000010) && ({row_reg, col_reg}<22'b0001001100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001100010000101101) && ({row_reg, col_reg}<22'b0001001100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001100100001010111) && ({row_reg, col_reg}<22'b0001001100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001100100010000010) && ({row_reg, col_reg}<22'b0001001100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001100100111010111) && ({row_reg, col_reg}<22'b0001001100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001001100101000000010) && ({row_reg, col_reg}<22'b0001001100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001100101010000010) && ({row_reg, col_reg}<22'b0001001100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001100101010101101) && ({row_reg, col_reg}<22'b0001001100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001100110000000010) && ({row_reg, col_reg}<22'b0001001100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001100110000101101) && ({row_reg, col_reg}<22'b0001001101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001101000001010111) && ({row_reg, col_reg}<22'b0001001101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001101000010000010) && ({row_reg, col_reg}<22'b0001001101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001101000111010111) && ({row_reg, col_reg}<22'b0001001101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001001101001000000010) && ({row_reg, col_reg}<22'b0001001101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001101001010000010) && ({row_reg, col_reg}<22'b0001001101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001101001010101101) && ({row_reg, col_reg}<22'b0001001101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001101010000000010) && ({row_reg, col_reg}<22'b0001001101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001101010000101101) && ({row_reg, col_reg}<22'b0001001101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001101100001010111) && ({row_reg, col_reg}<22'b0001001101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001101100010000010) && ({row_reg, col_reg}<22'b0001001101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001101100111010111) && ({row_reg, col_reg}<22'b0001001101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001001101101000000010) && ({row_reg, col_reg}<22'b0001001101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001101101010000010) && ({row_reg, col_reg}<22'b0001001101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001101101010101101) && ({row_reg, col_reg}<22'b0001001101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001101110000000010) && ({row_reg, col_reg}<22'b0001001101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001101110000101101) && ({row_reg, col_reg}<22'b0001001110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001110000001010111) && ({row_reg, col_reg}<22'b0001001110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001001110000010000010) && ({row_reg, col_reg}<22'b0001001110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001110000111010111) && ({row_reg, col_reg}<22'b0001001110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001001110001000000010) && ({row_reg, col_reg}<22'b0001001110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001110001010000010) && ({row_reg, col_reg}<22'b0001001110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001110001010101101) && ({row_reg, col_reg}<22'b0001001110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001110010000000010) && ({row_reg, col_reg}<22'b0001001110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001110010000101101) && ({row_reg, col_reg}<22'b0001001110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001110100001010111) && ({row_reg, col_reg}<22'b0001001110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001001110100010000010) && ({row_reg, col_reg}<22'b0001001110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001110100111010111) && ({row_reg, col_reg}<22'b0001001110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001001110101000000010) && ({row_reg, col_reg}<22'b0001001110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001110101010000010) && ({row_reg, col_reg}<22'b0001001110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001110101010101101) && ({row_reg, col_reg}<22'b0001001110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001110110000000010) && ({row_reg, col_reg}<22'b0001001110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001110110000101101) && ({row_reg, col_reg}<22'b0001001111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001111000001010111) && ({row_reg, col_reg}<22'b0001001111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001001111000010000010) && ({row_reg, col_reg}<22'b0001001111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001111000111010111) && ({row_reg, col_reg}<22'b0001001111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001001111001000000010) && ({row_reg, col_reg}<22'b0001001111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001111001010000010) && ({row_reg, col_reg}<22'b0001001111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001111001010101101) && ({row_reg, col_reg}<22'b0001001111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001111010000000010) && ({row_reg, col_reg}<22'b0001001111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001111010000101101) && ({row_reg, col_reg}<22'b0001001111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001111100001010111) && ({row_reg, col_reg}<22'b0001001111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001001111100010000010) && ({row_reg, col_reg}<22'b0001001111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001001111100111010111) && ({row_reg, col_reg}<22'b0001001111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001001111101000000010) && ({row_reg, col_reg}<22'b0001001111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001111101010000010) && ({row_reg, col_reg}<22'b0001001111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001111101010101101) && ({row_reg, col_reg}<22'b0001001111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001001111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001001111110000000010) && ({row_reg, col_reg}<22'b0001001111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001001111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001001111110000101101) && ({row_reg, col_reg}<22'b0001010000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010000000001010111) && ({row_reg, col_reg}<22'b0001010000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001010000000010000010) && ({row_reg, col_reg}<22'b0001010000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010000000111010111) && ({row_reg, col_reg}<22'b0001010000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010000001000000010) && ({row_reg, col_reg}<22'b0001010000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010000001010000010) && ({row_reg, col_reg}<22'b0001010000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010000001010101101) && ({row_reg, col_reg}<22'b0001010000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010000010000000010) && ({row_reg, col_reg}<22'b0001010000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010000010000101101) && ({row_reg, col_reg}<22'b0001010000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010000100001010111) && ({row_reg, col_reg}<22'b0001010000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001010000100010000010) && ({row_reg, col_reg}<22'b0001010000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010000100111010111) && ({row_reg, col_reg}<22'b0001010000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010000101000000010) && ({row_reg, col_reg}<22'b0001010000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010000101010000010) && ({row_reg, col_reg}<22'b0001010000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010000101010101101) && ({row_reg, col_reg}<22'b0001010000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010000110000000010) && ({row_reg, col_reg}<22'b0001010000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010000110000101101) && ({row_reg, col_reg}<22'b0001010001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010001000001010111) && ({row_reg, col_reg}<22'b0001010001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001010001000010000010) && ({row_reg, col_reg}<22'b0001010001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010001000111010111) && ({row_reg, col_reg}<22'b0001010001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010001001000000010) && ({row_reg, col_reg}<22'b0001010001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010001001010000010) && ({row_reg, col_reg}<22'b0001010001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010001001010101101) && ({row_reg, col_reg}<22'b0001010001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010001010000000010) && ({row_reg, col_reg}<22'b0001010001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010001010000101101) && ({row_reg, col_reg}<22'b0001010001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010001100001010111) && ({row_reg, col_reg}<22'b0001010001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010001100010000010) && ({row_reg, col_reg}<22'b0001010001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010001100111010111) && ({row_reg, col_reg}<22'b0001010001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010001101000000010) && ({row_reg, col_reg}<22'b0001010001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010001101010000010) && ({row_reg, col_reg}<22'b0001010001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010001101010101101) && ({row_reg, col_reg}<22'b0001010001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010001110000000010) && ({row_reg, col_reg}<22'b0001010001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010001110000101101) && ({row_reg, col_reg}<22'b0001010010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010010000001010111) && ({row_reg, col_reg}<22'b0001010010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010010000010000010) && ({row_reg, col_reg}<22'b0001010010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010010000111010111) && ({row_reg, col_reg}<22'b0001010010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010010001000000010) && ({row_reg, col_reg}<22'b0001010010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010010001010000010) && ({row_reg, col_reg}<22'b0001010010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010010001010101101) && ({row_reg, col_reg}<22'b0001010010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010010010000000010) && ({row_reg, col_reg}<22'b0001010010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010010010000101101) && ({row_reg, col_reg}<22'b0001010010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010010100001010111) && ({row_reg, col_reg}<22'b0001010010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010010100010000010) && ({row_reg, col_reg}<22'b0001010010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010010100111010111) && ({row_reg, col_reg}<22'b0001010010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010010101000000010) && ({row_reg, col_reg}<22'b0001010010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010010101010000010) && ({row_reg, col_reg}<22'b0001010010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010010101010101101) && ({row_reg, col_reg}<22'b0001010010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010010110000000010) && ({row_reg, col_reg}<22'b0001010010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010010110000101101) && ({row_reg, col_reg}<22'b0001010011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010011000001010111) && ({row_reg, col_reg}<22'b0001010011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010011000010000010) && ({row_reg, col_reg}<22'b0001010011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010011000111010111) && ({row_reg, col_reg}<22'b0001010011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010011001000000010) && ({row_reg, col_reg}<22'b0001010011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010011001010000010) && ({row_reg, col_reg}<22'b0001010011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010011001010101101) && ({row_reg, col_reg}<22'b0001010011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010011010000000010) && ({row_reg, col_reg}<22'b0001010011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010011010000101101) && ({row_reg, col_reg}<22'b0001010011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010011100001010111) && ({row_reg, col_reg}<22'b0001010011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010011100010000010) && ({row_reg, col_reg}<22'b0001010011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010011100111010111) && ({row_reg, col_reg}<22'b0001010011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010011101000000010) && ({row_reg, col_reg}<22'b0001010011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010011101010000010) && ({row_reg, col_reg}<22'b0001010011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010011101010101101) && ({row_reg, col_reg}<22'b0001010011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010011110000000010) && ({row_reg, col_reg}<22'b0001010011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010011110000101101) && ({row_reg, col_reg}<22'b0001010100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010100000001010111) && ({row_reg, col_reg}<22'b0001010100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010100000010000010) && ({row_reg, col_reg}<22'b0001010100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010100000111010111) && ({row_reg, col_reg}<22'b0001010100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010100001000000010) && ({row_reg, col_reg}<22'b0001010100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010100001010000010) && ({row_reg, col_reg}<22'b0001010100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010100001010101101) && ({row_reg, col_reg}<22'b0001010100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010100010000000010) && ({row_reg, col_reg}<22'b0001010100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010100010000101101) && ({row_reg, col_reg}<22'b0001010100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010100100001010111) && ({row_reg, col_reg}<22'b0001010100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010100100010000010) && ({row_reg, col_reg}<22'b0001010100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010100100111010111) && ({row_reg, col_reg}<22'b0001010100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010100101000000010) && ({row_reg, col_reg}<22'b0001010100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010100101010000010) && ({row_reg, col_reg}<22'b0001010100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010100101010101101) && ({row_reg, col_reg}<22'b0001010100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010100110000000010) && ({row_reg, col_reg}<22'b0001010100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010100110000101101) && ({row_reg, col_reg}<22'b0001010101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010101000001010111) && ({row_reg, col_reg}<22'b0001010101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010101000010000010) && ({row_reg, col_reg}<22'b0001010101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010101000111010111) && ({row_reg, col_reg}<22'b0001010101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010101001000000010) && ({row_reg, col_reg}<22'b0001010101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010101001010000010) && ({row_reg, col_reg}<22'b0001010101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010101001010101101) && ({row_reg, col_reg}<22'b0001010101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010101010000000010) && ({row_reg, col_reg}<22'b0001010101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010101010000101101) && ({row_reg, col_reg}<22'b0001010101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010101100001010111) && ({row_reg, col_reg}<22'b0001010101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010101100010000010) && ({row_reg, col_reg}<22'b0001010101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010101100111010111) && ({row_reg, col_reg}<22'b0001010101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010101101000000010) && ({row_reg, col_reg}<22'b0001010101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010101101010000010) && ({row_reg, col_reg}<22'b0001010101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010101101010101101) && ({row_reg, col_reg}<22'b0001010101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010101110000000010) && ({row_reg, col_reg}<22'b0001010101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010101110000101101) && ({row_reg, col_reg}<22'b0001010110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010110000001010111) && ({row_reg, col_reg}<22'b0001010110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010110000010000010) && ({row_reg, col_reg}<22'b0001010110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010110000111010111) && ({row_reg, col_reg}<22'b0001010110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001010110001000000010) && ({row_reg, col_reg}<22'b0001010110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010110001010000010) && ({row_reg, col_reg}<22'b0001010110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010110001010101101) && ({row_reg, col_reg}<22'b0001010110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010110010000000010) && ({row_reg, col_reg}<22'b0001010110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010110010000101101) && ({row_reg, col_reg}<22'b0001010110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010110100001010111) && ({row_reg, col_reg}<22'b0001010110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010110100010000010) && ({row_reg, col_reg}<22'b0001010110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010110100111010111) && ({row_reg, col_reg}<22'b0001010110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001010110101000000010) && ({row_reg, col_reg}<22'b0001010110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010110101010000010) && ({row_reg, col_reg}<22'b0001010110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010110101010101101) && ({row_reg, col_reg}<22'b0001010110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010110110000000010) && ({row_reg, col_reg}<22'b0001010110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010110110000101101) && ({row_reg, col_reg}<22'b0001010111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010111000001010111) && ({row_reg, col_reg}<22'b0001010111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010111000010000010) && ({row_reg, col_reg}<22'b0001010111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010111000111010111) && ({row_reg, col_reg}<22'b0001010111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001010111001000000010) && ({row_reg, col_reg}<22'b0001010111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010111001010000010) && ({row_reg, col_reg}<22'b0001010111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010111001010101101) && ({row_reg, col_reg}<22'b0001010111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010111010000000010) && ({row_reg, col_reg}<22'b0001010111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010111010000101101) && ({row_reg, col_reg}<22'b0001010111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010111100001010111) && ({row_reg, col_reg}<22'b0001010111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001010111100010000010) && ({row_reg, col_reg}<22'b0001010111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001010111100111010111) && ({row_reg, col_reg}<22'b0001010111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001010111101000000010) && ({row_reg, col_reg}<22'b0001010111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010111101010000010) && ({row_reg, col_reg}<22'b0001010111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010111101010101101) && ({row_reg, col_reg}<22'b0001010111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001010111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001010111110000000010) && ({row_reg, col_reg}<22'b0001010111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001010111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001010111110000101101) && ({row_reg, col_reg}<22'b0001011000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011000000001010111) && ({row_reg, col_reg}<22'b0001011000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001011000000010000010) && ({row_reg, col_reg}<22'b0001011000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011000000111010111) && ({row_reg, col_reg}<22'b0001011000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001011000001000000010) && ({row_reg, col_reg}<22'b0001011000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011000001010000010) && ({row_reg, col_reg}<22'b0001011000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011000001010101101) && ({row_reg, col_reg}<22'b0001011000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011000010000000010) && ({row_reg, col_reg}<22'b0001011000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011000010000101101) && ({row_reg, col_reg}<22'b0001011000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011000100001010111) && ({row_reg, col_reg}<22'b0001011000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001011000100010000010) && ({row_reg, col_reg}<22'b0001011000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011000100111010111) && ({row_reg, col_reg}<22'b0001011000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001011000101000000010) && ({row_reg, col_reg}<22'b0001011000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011000101010000010) && ({row_reg, col_reg}<22'b0001011000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011000101010101101) && ({row_reg, col_reg}<22'b0001011000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011000110000000010) && ({row_reg, col_reg}<22'b0001011000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011000110000101101) && ({row_reg, col_reg}<22'b0001011001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011001000001010111) && ({row_reg, col_reg}<22'b0001011001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001011001000010000010) && ({row_reg, col_reg}<22'b0001011001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011001000111010111) && ({row_reg, col_reg}<22'b0001011001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001011001001000000010) && ({row_reg, col_reg}<22'b0001011001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011001001010000010) && ({row_reg, col_reg}<22'b0001011001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011001001010101101) && ({row_reg, col_reg}<22'b0001011001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011001010000000010) && ({row_reg, col_reg}<22'b0001011001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011001010000101101) && ({row_reg, col_reg}<22'b0001011001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011001100001010111) && ({row_reg, col_reg}<22'b0001011001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001011001100010000010) && ({row_reg, col_reg}<22'b0001011001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011001100111010111) && ({row_reg, col_reg}<22'b0001011001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011001101000000010) && ({row_reg, col_reg}<22'b0001011001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011001101010000010) && ({row_reg, col_reg}<22'b0001011001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011001101010101101) && ({row_reg, col_reg}<22'b0001011001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011001110000000010) && ({row_reg, col_reg}<22'b0001011001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011001110000101101) && ({row_reg, col_reg}<22'b0001011010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011010000001010111) && ({row_reg, col_reg}<22'b0001011010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001011010000010000010) && ({row_reg, col_reg}<22'b0001011010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011010000111010111) && ({row_reg, col_reg}<22'b0001011010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011010001000000010) && ({row_reg, col_reg}<22'b0001011010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011010001010000010) && ({row_reg, col_reg}<22'b0001011010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011010001010101101) && ({row_reg, col_reg}<22'b0001011010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011010010000000010) && ({row_reg, col_reg}<22'b0001011010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011010010000101101) && ({row_reg, col_reg}<22'b0001011010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011010100001010111) && ({row_reg, col_reg}<22'b0001011010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001011010100010000010) && ({row_reg, col_reg}<22'b0001011010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011010100111010111) && ({row_reg, col_reg}<22'b0001011010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011010101000000010) && ({row_reg, col_reg}<22'b0001011010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011010101010000010) && ({row_reg, col_reg}<22'b0001011010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011010101010101101) && ({row_reg, col_reg}<22'b0001011010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011010110000000010) && ({row_reg, col_reg}<22'b0001011010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011010110000101101) && ({row_reg, col_reg}<22'b0001011011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011011000001010111) && ({row_reg, col_reg}<22'b0001011011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001011011000010000010) && ({row_reg, col_reg}<22'b0001011011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011011000111010111) && ({row_reg, col_reg}<22'b0001011011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011011001000000010) && ({row_reg, col_reg}<22'b0001011011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011011001010000010) && ({row_reg, col_reg}<22'b0001011011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011011001010101101) && ({row_reg, col_reg}<22'b0001011011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011011010000000010) && ({row_reg, col_reg}<22'b0001011011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011011010000101101) && ({row_reg, col_reg}<22'b0001011011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011011100001010111) && ({row_reg, col_reg}<22'b0001011011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011011100010000010) && ({row_reg, col_reg}<22'b0001011011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011011100111010111) && ({row_reg, col_reg}<22'b0001011011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011011101000000010) && ({row_reg, col_reg}<22'b0001011011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011011101010000010) && ({row_reg, col_reg}<22'b0001011011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011011101010101101) && ({row_reg, col_reg}<22'b0001011011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011011110000000010) && ({row_reg, col_reg}<22'b0001011011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011011110000101101) && ({row_reg, col_reg}<22'b0001011100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011100000001010111) && ({row_reg, col_reg}<22'b0001011100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011100000010000010) && ({row_reg, col_reg}<22'b0001011100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011100000111010111) && ({row_reg, col_reg}<22'b0001011100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011100001000000010) && ({row_reg, col_reg}<22'b0001011100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011100001010000010) && ({row_reg, col_reg}<22'b0001011100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011100001010101101) && ({row_reg, col_reg}<22'b0001011100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011100010000000010) && ({row_reg, col_reg}<22'b0001011100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011100010000101101) && ({row_reg, col_reg}<22'b0001011100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011100100001010111) && ({row_reg, col_reg}<22'b0001011100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011100100010000010) && ({row_reg, col_reg}<22'b0001011100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011100100111010111) && ({row_reg, col_reg}<22'b0001011100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011100101000000010) && ({row_reg, col_reg}<22'b0001011100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011100101010000010) && ({row_reg, col_reg}<22'b0001011100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011100101010101101) && ({row_reg, col_reg}<22'b0001011100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011100110000000010) && ({row_reg, col_reg}<22'b0001011100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011100110000101101) && ({row_reg, col_reg}<22'b0001011101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011101000001010111) && ({row_reg, col_reg}<22'b0001011101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011101000010000010) && ({row_reg, col_reg}<22'b0001011101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011101000111010111) && ({row_reg, col_reg}<22'b0001011101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011101001000000010) && ({row_reg, col_reg}<22'b0001011101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011101001010000010) && ({row_reg, col_reg}<22'b0001011101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011101001010101101) && ({row_reg, col_reg}<22'b0001011101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011101010000000010) && ({row_reg, col_reg}<22'b0001011101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011101010000101101) && ({row_reg, col_reg}<22'b0001011101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011101100001010111) && ({row_reg, col_reg}<22'b0001011101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011101100010000010) && ({row_reg, col_reg}<22'b0001011101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011101100111010111) && ({row_reg, col_reg}<22'b0001011101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011101101000000010) && ({row_reg, col_reg}<22'b0001011101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011101101010000010) && ({row_reg, col_reg}<22'b0001011101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011101101010101101) && ({row_reg, col_reg}<22'b0001011101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011101110000000010) && ({row_reg, col_reg}<22'b0001011101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011101110000101101) && ({row_reg, col_reg}<22'b0001011110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011110000001010111) && ({row_reg, col_reg}<22'b0001011110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011110000010000010) && ({row_reg, col_reg}<22'b0001011110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011110000111010111) && ({row_reg, col_reg}<22'b0001011110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011110001000000010) && ({row_reg, col_reg}<22'b0001011110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011110001010000010) && ({row_reg, col_reg}<22'b0001011110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011110001010101101) && ({row_reg, col_reg}<22'b0001011110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011110010000000010) && ({row_reg, col_reg}<22'b0001011110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011110010000101101) && ({row_reg, col_reg}<22'b0001011110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011110100001010111) && ({row_reg, col_reg}<22'b0001011110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011110100010000010) && ({row_reg, col_reg}<22'b0001011110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011110100111010111) && ({row_reg, col_reg}<22'b0001011110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011110101000000010) && ({row_reg, col_reg}<22'b0001011110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011110101010000010) && ({row_reg, col_reg}<22'b0001011110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011110101010101101) && ({row_reg, col_reg}<22'b0001011110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011110110000000010) && ({row_reg, col_reg}<22'b0001011110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011110110000101101) && ({row_reg, col_reg}<22'b0001011111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011111000001010111) && ({row_reg, col_reg}<22'b0001011111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011111000010000010) && ({row_reg, col_reg}<22'b0001011111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011111000111010111) && ({row_reg, col_reg}<22'b0001011111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011111001000000010) && ({row_reg, col_reg}<22'b0001011111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011111001010000010) && ({row_reg, col_reg}<22'b0001011111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011111001010101101) && ({row_reg, col_reg}<22'b0001011111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011111010000000010) && ({row_reg, col_reg}<22'b0001011111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011111010000101101) && ({row_reg, col_reg}<22'b0001011111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011111100001010111) && ({row_reg, col_reg}<22'b0001011111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011111100010000010) && ({row_reg, col_reg}<22'b0001011111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001011111100111010111) && ({row_reg, col_reg}<22'b0001011111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001011111101000000010) && ({row_reg, col_reg}<22'b0001011111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011111101010000010) && ({row_reg, col_reg}<22'b0001011111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011111101010101101) && ({row_reg, col_reg}<22'b0001011111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001011111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001011111110000000010) && ({row_reg, col_reg}<22'b0001011111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001011111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001011111110000101101) && ({row_reg, col_reg}<22'b0001100000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100000000001010111) && ({row_reg, col_reg}<22'b0001100000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100000000010000010) && ({row_reg, col_reg}<22'b0001100000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100000000111010111) && ({row_reg, col_reg}<22'b0001100000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100000001000000010) && ({row_reg, col_reg}<22'b0001100000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100000001010000010) && ({row_reg, col_reg}<22'b0001100000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100000001010101101) && ({row_reg, col_reg}<22'b0001100000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100000010000000010) && ({row_reg, col_reg}<22'b0001100000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100000010000101101) && ({row_reg, col_reg}<22'b0001100000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100000100001010111) && ({row_reg, col_reg}<22'b0001100000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100000100010000010) && ({row_reg, col_reg}<22'b0001100000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100000100111010111) && ({row_reg, col_reg}<22'b0001100000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100000101000000010) && ({row_reg, col_reg}<22'b0001100000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100000101010000010) && ({row_reg, col_reg}<22'b0001100000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100000101010101101) && ({row_reg, col_reg}<22'b0001100000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100000110000000010) && ({row_reg, col_reg}<22'b0001100000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100000110000101101) && ({row_reg, col_reg}<22'b0001100001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100001000001010111) && ({row_reg, col_reg}<22'b0001100001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100001000010000010) && ({row_reg, col_reg}<22'b0001100001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100001000111010111) && ({row_reg, col_reg}<22'b0001100001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001100001001000000010) && ({row_reg, col_reg}<22'b0001100001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100001001010000010) && ({row_reg, col_reg}<22'b0001100001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100001001010101101) && ({row_reg, col_reg}<22'b0001100001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100001010000000010) && ({row_reg, col_reg}<22'b0001100001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100001010000101101) && ({row_reg, col_reg}<22'b0001100001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100001100001010111) && ({row_reg, col_reg}<22'b0001100001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100001100010000010) && ({row_reg, col_reg}<22'b0001100001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100001100111010111) && ({row_reg, col_reg}<22'b0001100001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001100001101000000010) && ({row_reg, col_reg}<22'b0001100001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100001101010000010) && ({row_reg, col_reg}<22'b0001100001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100001101010101101) && ({row_reg, col_reg}<22'b0001100001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100001110000000010) && ({row_reg, col_reg}<22'b0001100001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100001110000101101) && ({row_reg, col_reg}<22'b0001100010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100010000001010111) && ({row_reg, col_reg}<22'b0001100010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100010000010000010) && ({row_reg, col_reg}<22'b0001100010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100010000111010111) && ({row_reg, col_reg}<22'b0001100010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001100010001000000010) && ({row_reg, col_reg}<22'b0001100010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100010001010000010) && ({row_reg, col_reg}<22'b0001100010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100010001010101101) && ({row_reg, col_reg}<22'b0001100010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100010010000000010) && ({row_reg, col_reg}<22'b0001100010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100010010000101101) && ({row_reg, col_reg}<22'b0001100010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100010100001010111) && ({row_reg, col_reg}<22'b0001100010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100010100010000010) && ({row_reg, col_reg}<22'b0001100010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100010100111010111) && ({row_reg, col_reg}<22'b0001100010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100010101000000010) && ({row_reg, col_reg}<22'b0001100010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100010101010000010) && ({row_reg, col_reg}<22'b0001100010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100010101010101101) && ({row_reg, col_reg}<22'b0001100010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100010110000000010) && ({row_reg, col_reg}<22'b0001100010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100010110000101101) && ({row_reg, col_reg}<22'b0001100011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100011000001010111) && ({row_reg, col_reg}<22'b0001100011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001100011000010000010) && ({row_reg, col_reg}<22'b0001100011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100011000111010111) && ({row_reg, col_reg}<22'b0001100011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100011001000000010) && ({row_reg, col_reg}<22'b0001100011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100011001010000010) && ({row_reg, col_reg}<22'b0001100011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100011001010101101) && ({row_reg, col_reg}<22'b0001100011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100011010000000010) && ({row_reg, col_reg}<22'b0001100011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100011010000101101) && ({row_reg, col_reg}<22'b0001100011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100011100001010111) && ({row_reg, col_reg}<22'b0001100011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001100011100010000010) && ({row_reg, col_reg}<22'b0001100011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100011100111010111) && ({row_reg, col_reg}<22'b0001100011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100011101000000010) && ({row_reg, col_reg}<22'b0001100011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100011101010000010) && ({row_reg, col_reg}<22'b0001100011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100011101010101101) && ({row_reg, col_reg}<22'b0001100011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100011110000000010) && ({row_reg, col_reg}<22'b0001100011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100011110000101101) && ({row_reg, col_reg}<22'b0001100100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100100000001010111) && ({row_reg, col_reg}<22'b0001100100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001100100000010000010) && ({row_reg, col_reg}<22'b0001100100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100100000111010111) && ({row_reg, col_reg}<22'b0001100100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100100001000000010) && ({row_reg, col_reg}<22'b0001100100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100100001010000010) && ({row_reg, col_reg}<22'b0001100100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100100001010101101) && ({row_reg, col_reg}<22'b0001100100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100100010000000010) && ({row_reg, col_reg}<22'b0001100100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100100010000101101) && ({row_reg, col_reg}<22'b0001100100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100100100001010111) && ({row_reg, col_reg}<22'b0001100100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100100100010000010) && ({row_reg, col_reg}<22'b0001100100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100100100111010111) && ({row_reg, col_reg}<22'b0001100100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100100101000000010) && ({row_reg, col_reg}<22'b0001100100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100100101010000010) && ({row_reg, col_reg}<22'b0001100100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100100101010101101) && ({row_reg, col_reg}<22'b0001100100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100100110000000010) && ({row_reg, col_reg}<22'b0001100100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100100110000101101) && ({row_reg, col_reg}<22'b0001100101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100101000001010111) && ({row_reg, col_reg}<22'b0001100101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001100101000010000010) && ({row_reg, col_reg}<22'b0001100101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100101000111010111) && ({row_reg, col_reg}<22'b0001100101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100101001000000010) && ({row_reg, col_reg}<22'b0001100101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100101001010000010) && ({row_reg, col_reg}<22'b0001100101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100101001010101101) && ({row_reg, col_reg}<22'b0001100101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100101010000000010) && ({row_reg, col_reg}<22'b0001100101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100101010000101101) && ({row_reg, col_reg}<22'b0001100101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100101100001010111) && ({row_reg, col_reg}<22'b0001100101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100101100010000010) && ({row_reg, col_reg}<22'b0001100101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100101100111010111) && ({row_reg, col_reg}<22'b0001100101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100101101000000010) && ({row_reg, col_reg}<22'b0001100101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100101101010000010) && ({row_reg, col_reg}<22'b0001100101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100101101010101101) && ({row_reg, col_reg}<22'b0001100101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100101110000000010) && ({row_reg, col_reg}<22'b0001100101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100101110000101101) && ({row_reg, col_reg}<22'b0001100110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100110000001010111) && ({row_reg, col_reg}<22'b0001100110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100110000010000010) && ({row_reg, col_reg}<22'b0001100110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100110000111010111) && ({row_reg, col_reg}<22'b0001100110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100110001000000010) && ({row_reg, col_reg}<22'b0001100110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100110001010000010) && ({row_reg, col_reg}<22'b0001100110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100110001010101101) && ({row_reg, col_reg}<22'b0001100110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100110010000000010) && ({row_reg, col_reg}<22'b0001100110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100110010000101101) && ({row_reg, col_reg}<22'b0001100110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100110100001010111) && ({row_reg, col_reg}<22'b0001100110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100110100010000010) && ({row_reg, col_reg}<22'b0001100110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100110100111010111) && ({row_reg, col_reg}<22'b0001100110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100110101000000010) && ({row_reg, col_reg}<22'b0001100110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100110101010000010) && ({row_reg, col_reg}<22'b0001100110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100110101010101101) && ({row_reg, col_reg}<22'b0001100110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100110110000000010) && ({row_reg, col_reg}<22'b0001100110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100110110000101101) && ({row_reg, col_reg}<22'b0001100111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100111000001010111) && ({row_reg, col_reg}<22'b0001100111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100111000010000010) && ({row_reg, col_reg}<22'b0001100111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100111000111010111) && ({row_reg, col_reg}<22'b0001100111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100111001000000010) && ({row_reg, col_reg}<22'b0001100111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100111001010000010) && ({row_reg, col_reg}<22'b0001100111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100111001010101101) && ({row_reg, col_reg}<22'b0001100111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100111010000000010) && ({row_reg, col_reg}<22'b0001100111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100111010000101101) && ({row_reg, col_reg}<22'b0001100111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100111100001010111) && ({row_reg, col_reg}<22'b0001100111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100111100010000010) && ({row_reg, col_reg}<22'b0001100111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001100111100111010111) && ({row_reg, col_reg}<22'b0001100111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001100111101000000010) && ({row_reg, col_reg}<22'b0001100111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100111101010000010) && ({row_reg, col_reg}<22'b0001100111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100111101010101101) && ({row_reg, col_reg}<22'b0001100111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001100111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001100111110000000010) && ({row_reg, col_reg}<22'b0001100111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001100111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001100111110000101101) && ({row_reg, col_reg}<22'b0001101000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101000000001010111) && ({row_reg, col_reg}<22'b0001101000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101000000010000010) && ({row_reg, col_reg}<22'b0001101000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101000000111010111) && ({row_reg, col_reg}<22'b0001101000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101000001000000010) && ({row_reg, col_reg}<22'b0001101000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101000001010000010) && ({row_reg, col_reg}<22'b0001101000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101000001010101101) && ({row_reg, col_reg}<22'b0001101000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101000010000000010) && ({row_reg, col_reg}<22'b0001101000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101000010000101101) && ({row_reg, col_reg}<22'b0001101000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101000100001010111) && ({row_reg, col_reg}<22'b0001101000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101000100010000010) && ({row_reg, col_reg}<22'b0001101000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101000100111010111) && ({row_reg, col_reg}<22'b0001101000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101000101000000010) && ({row_reg, col_reg}<22'b0001101000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101000101010000010) && ({row_reg, col_reg}<22'b0001101000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101000101010101101) && ({row_reg, col_reg}<22'b0001101000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101000110000000010) && ({row_reg, col_reg}<22'b0001101000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101000110000101101) && ({row_reg, col_reg}<22'b0001101001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101001000001010111) && ({row_reg, col_reg}<22'b0001101001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101001000010000010) && ({row_reg, col_reg}<22'b0001101001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101001000111010111) && ({row_reg, col_reg}<22'b0001101001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101001001000000010) && ({row_reg, col_reg}<22'b0001101001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101001001010000010) && ({row_reg, col_reg}<22'b0001101001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101001001010101101) && ({row_reg, col_reg}<22'b0001101001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101001010000000010) && ({row_reg, col_reg}<22'b0001101001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101001010000101101) && ({row_reg, col_reg}<22'b0001101001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101001100001010111) && ({row_reg, col_reg}<22'b0001101001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101001100010000010) && ({row_reg, col_reg}<22'b0001101001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101001100111010111) && ({row_reg, col_reg}<22'b0001101001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101001101000000010) && ({row_reg, col_reg}<22'b0001101001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101001101010000010) && ({row_reg, col_reg}<22'b0001101001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101001101010101101) && ({row_reg, col_reg}<22'b0001101001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101001110000000010) && ({row_reg, col_reg}<22'b0001101001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101001110000101101) && ({row_reg, col_reg}<22'b0001101010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101010000001010111) && ({row_reg, col_reg}<22'b0001101010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101010000010000010) && ({row_reg, col_reg}<22'b0001101010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101010000111010111) && ({row_reg, col_reg}<22'b0001101010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101010001000000010) && ({row_reg, col_reg}<22'b0001101010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101010001010000010) && ({row_reg, col_reg}<22'b0001101010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101010001010101101) && ({row_reg, col_reg}<22'b0001101010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101010010000000010) && ({row_reg, col_reg}<22'b0001101010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101010010000101101) && ({row_reg, col_reg}<22'b0001101010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101010100001010111) && ({row_reg, col_reg}<22'b0001101010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101010100010000010) && ({row_reg, col_reg}<22'b0001101010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101010100111010111) && ({row_reg, col_reg}<22'b0001101010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101010101000000010) && ({row_reg, col_reg}<22'b0001101010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101010101010000010) && ({row_reg, col_reg}<22'b0001101010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101010101010101101) && ({row_reg, col_reg}<22'b0001101010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101010110000000010) && ({row_reg, col_reg}<22'b0001101010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101010110000101101) && ({row_reg, col_reg}<22'b0001101011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101011000001010111) && ({row_reg, col_reg}<22'b0001101011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101011000010000010) && ({row_reg, col_reg}<22'b0001101011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101011000111010111) && ({row_reg, col_reg}<22'b0001101011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001101011001000000010) && ({row_reg, col_reg}<22'b0001101011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101011001010000010) && ({row_reg, col_reg}<22'b0001101011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101011001010101101) && ({row_reg, col_reg}<22'b0001101011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101011010000000010) && ({row_reg, col_reg}<22'b0001101011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101011010000101101) && ({row_reg, col_reg}<22'b0001101011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101011100001010111) && ({row_reg, col_reg}<22'b0001101011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101011100010000010) && ({row_reg, col_reg}<22'b0001101011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101011100111010111) && ({row_reg, col_reg}<22'b0001101011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001101011101000000010) && ({row_reg, col_reg}<22'b0001101011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101011101010000010) && ({row_reg, col_reg}<22'b0001101011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101011101010101101) && ({row_reg, col_reg}<22'b0001101011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101011110000000010) && ({row_reg, col_reg}<22'b0001101011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101011110000101101) && ({row_reg, col_reg}<22'b0001101100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101100000001010111) && ({row_reg, col_reg}<22'b0001101100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101100000010000010) && ({row_reg, col_reg}<22'b0001101100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101100000111010111) && ({row_reg, col_reg}<22'b0001101100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001101100001000000010) && ({row_reg, col_reg}<22'b0001101100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101100001010000010) && ({row_reg, col_reg}<22'b0001101100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101100001010101101) && ({row_reg, col_reg}<22'b0001101100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101100010000000010) && ({row_reg, col_reg}<22'b0001101100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101100010000101101) && ({row_reg, col_reg}<22'b0001101100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101100100001010111) && ({row_reg, col_reg}<22'b0001101100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101100100010000010) && ({row_reg, col_reg}<22'b0001101100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101100100111010111) && ({row_reg, col_reg}<22'b0001101100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101100101000000010) && ({row_reg, col_reg}<22'b0001101100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101100101010000010) && ({row_reg, col_reg}<22'b0001101100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101100101010101101) && ({row_reg, col_reg}<22'b0001101100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101100110000000010) && ({row_reg, col_reg}<22'b0001101100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101100110000101101) && ({row_reg, col_reg}<22'b0001101101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101101000001010111) && ({row_reg, col_reg}<22'b0001101101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001101101000010000010) && ({row_reg, col_reg}<22'b0001101101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101101000111010111) && ({row_reg, col_reg}<22'b0001101101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101101001000000010) && ({row_reg, col_reg}<22'b0001101101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101101001010000010) && ({row_reg, col_reg}<22'b0001101101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101101001010101101) && ({row_reg, col_reg}<22'b0001101101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101101010000000010) && ({row_reg, col_reg}<22'b0001101101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101101010000101101) && ({row_reg, col_reg}<22'b0001101101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101101100001010111) && ({row_reg, col_reg}<22'b0001101101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001101101100010000010) && ({row_reg, col_reg}<22'b0001101101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101101100111010111) && ({row_reg, col_reg}<22'b0001101101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101101101000000010) && ({row_reg, col_reg}<22'b0001101101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101101101010000010) && ({row_reg, col_reg}<22'b0001101101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101101101010101101) && ({row_reg, col_reg}<22'b0001101101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101101110000000010) && ({row_reg, col_reg}<22'b0001101101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101101110000101101) && ({row_reg, col_reg}<22'b0001101110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101110000001010111) && ({row_reg, col_reg}<22'b0001101110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001101110000010000010) && ({row_reg, col_reg}<22'b0001101110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101110000111010111) && ({row_reg, col_reg}<22'b0001101110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101110001000000010) && ({row_reg, col_reg}<22'b0001101110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101110001010000010) && ({row_reg, col_reg}<22'b0001101110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101110001010101101) && ({row_reg, col_reg}<22'b0001101110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101110010000000010) && ({row_reg, col_reg}<22'b0001101110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101110010000101101) && ({row_reg, col_reg}<22'b0001101110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101110100001010111) && ({row_reg, col_reg}<22'b0001101110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101110100010000010) && ({row_reg, col_reg}<22'b0001101110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101110100111010111) && ({row_reg, col_reg}<22'b0001101110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101110101000000010) && ({row_reg, col_reg}<22'b0001101110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101110101010000010) && ({row_reg, col_reg}<22'b0001101110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101110101010101101) && ({row_reg, col_reg}<22'b0001101110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101110110000000010) && ({row_reg, col_reg}<22'b0001101110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101110110000101101) && ({row_reg, col_reg}<22'b0001101111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101111000001010111) && ({row_reg, col_reg}<22'b0001101111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001101111000010000010) && ({row_reg, col_reg}<22'b0001101111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101111000111010111) && ({row_reg, col_reg}<22'b0001101111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101111001000000010) && ({row_reg, col_reg}<22'b0001101111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101111001010000010) && ({row_reg, col_reg}<22'b0001101111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101111001010101101) && ({row_reg, col_reg}<22'b0001101111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101111010000000010) && ({row_reg, col_reg}<22'b0001101111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101111010000101101) && ({row_reg, col_reg}<22'b0001101111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101111100001010111) && ({row_reg, col_reg}<22'b0001101111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101111100010000010) && ({row_reg, col_reg}<22'b0001101111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001101111100111010111) && ({row_reg, col_reg}<22'b0001101111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001101111101000000010) && ({row_reg, col_reg}<22'b0001101111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101111101010000010) && ({row_reg, col_reg}<22'b0001101111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101111101010101101) && ({row_reg, col_reg}<22'b0001101111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001101111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001101111110000000010) && ({row_reg, col_reg}<22'b0001101111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001101111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001101111110000101101) && ({row_reg, col_reg}<22'b0001110000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110000000001010111) && ({row_reg, col_reg}<22'b0001110000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110000000010000010) && ({row_reg, col_reg}<22'b0001110000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110000000111010111) && ({row_reg, col_reg}<22'b0001110000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110000001000000010) && ({row_reg, col_reg}<22'b0001110000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110000001010000010) && ({row_reg, col_reg}<22'b0001110000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110000001010101101) && ({row_reg, col_reg}<22'b0001110000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110000010000000010) && ({row_reg, col_reg}<22'b0001110000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110000010000101101) && ({row_reg, col_reg}<22'b0001110000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110000100001010111) && ({row_reg, col_reg}<22'b0001110000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110000100010000010) && ({row_reg, col_reg}<22'b0001110000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110000100111010111) && ({row_reg, col_reg}<22'b0001110000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110000101000000010) && ({row_reg, col_reg}<22'b0001110000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110000101010000010) && ({row_reg, col_reg}<22'b0001110000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110000101010101101) && ({row_reg, col_reg}<22'b0001110000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110000110000000010) && ({row_reg, col_reg}<22'b0001110000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110000110000101101) && ({row_reg, col_reg}<22'b0001110001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110001000001010111) && ({row_reg, col_reg}<22'b0001110001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110001000010000010) && ({row_reg, col_reg}<22'b0001110001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110001000111010111) && ({row_reg, col_reg}<22'b0001110001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110001001000000010) && ({row_reg, col_reg}<22'b0001110001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110001001010000010) && ({row_reg, col_reg}<22'b0001110001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110001001010101101) && ({row_reg, col_reg}<22'b0001110001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110001010000000010) && ({row_reg, col_reg}<22'b0001110001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110001010000101101) && ({row_reg, col_reg}<22'b0001110001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110001100001010111) && ({row_reg, col_reg}<22'b0001110001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110001100010000010) && ({row_reg, col_reg}<22'b0001110001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110001100111010111) && ({row_reg, col_reg}<22'b0001110001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110001101000000010) && ({row_reg, col_reg}<22'b0001110001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110001101010000010) && ({row_reg, col_reg}<22'b0001110001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110001101010101101) && ({row_reg, col_reg}<22'b0001110001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110001110000000010) && ({row_reg, col_reg}<22'b0001110001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110001110000101101) && ({row_reg, col_reg}<22'b0001110010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110010000001010111) && ({row_reg, col_reg}<22'b0001110010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110010000010000010) && ({row_reg, col_reg}<22'b0001110010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110010000111010111) && ({row_reg, col_reg}<22'b0001110010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110010001000000010) && ({row_reg, col_reg}<22'b0001110010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110010001010000010) && ({row_reg, col_reg}<22'b0001110010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110010001010101101) && ({row_reg, col_reg}<22'b0001110010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110010010000000010) && ({row_reg, col_reg}<22'b0001110010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110010010000101101) && ({row_reg, col_reg}<22'b0001110010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110010100001010111) && ({row_reg, col_reg}<22'b0001110010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110010100010000010) && ({row_reg, col_reg}<22'b0001110010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110010100111010111) && ({row_reg, col_reg}<22'b0001110010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110010101000000010) && ({row_reg, col_reg}<22'b0001110010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110010101010000010) && ({row_reg, col_reg}<22'b0001110010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110010101010101101) && ({row_reg, col_reg}<22'b0001110010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110010110000000010) && ({row_reg, col_reg}<22'b0001110010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110010110000101101) && ({row_reg, col_reg}<22'b0001110011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110011000001010111) && ({row_reg, col_reg}<22'b0001110011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110011000010000010) && ({row_reg, col_reg}<22'b0001110011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110011000111010111) && ({row_reg, col_reg}<22'b0001110011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110011001000000010) && ({row_reg, col_reg}<22'b0001110011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110011001010000010) && ({row_reg, col_reg}<22'b0001110011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110011001010101101) && ({row_reg, col_reg}<22'b0001110011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110011010000000010) && ({row_reg, col_reg}<22'b0001110011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110011010000101101) && ({row_reg, col_reg}<22'b0001110011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110011100001010111) && ({row_reg, col_reg}<22'b0001110011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110011100010000010) && ({row_reg, col_reg}<22'b0001110011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110011100111010111) && ({row_reg, col_reg}<22'b0001110011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110011101000000010) && ({row_reg, col_reg}<22'b0001110011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110011101010000010) && ({row_reg, col_reg}<22'b0001110011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110011101010101101) && ({row_reg, col_reg}<22'b0001110011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110011110000000010) && ({row_reg, col_reg}<22'b0001110011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110011110000101101) && ({row_reg, col_reg}<22'b0001110100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110100000001010111) && ({row_reg, col_reg}<22'b0001110100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110100000010000010) && ({row_reg, col_reg}<22'b0001110100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110100000111010111) && ({row_reg, col_reg}<22'b0001110100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001110100001000000010) && ({row_reg, col_reg}<22'b0001110100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110100001010000010) && ({row_reg, col_reg}<22'b0001110100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110100001010101101) && ({row_reg, col_reg}<22'b0001110100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110100010000000010) && ({row_reg, col_reg}<22'b0001110100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110100010000101101) && ({row_reg, col_reg}<22'b0001110100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110100100001010111) && ({row_reg, col_reg}<22'b0001110100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110100100010000010) && ({row_reg, col_reg}<22'b0001110100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110100100111010111) && ({row_reg, col_reg}<22'b0001110100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001110100101000000010) && ({row_reg, col_reg}<22'b0001110100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110100101010000010) && ({row_reg, col_reg}<22'b0001110100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110100101010101101) && ({row_reg, col_reg}<22'b0001110100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110100110000000010) && ({row_reg, col_reg}<22'b0001110100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110100110000101101) && ({row_reg, col_reg}<22'b0001110101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110101000001010111) && ({row_reg, col_reg}<22'b0001110101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101000010000010) && ({row_reg, col_reg}<22'b0001110101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110101000111010111) && ({row_reg, col_reg}<22'b0001110101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101001000000010) && ({row_reg, col_reg}<22'b0001110101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110101001010000010) && ({row_reg, col_reg}<22'b0001110101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110101001010101101) && ({row_reg, col_reg}<22'b0001110101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110101010000000010) && ({row_reg, col_reg}<22'b0001110101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110101010000101101) && ({row_reg, col_reg}<22'b0001110101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110101100001010111) && ({row_reg, col_reg}<22'b0001110101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100010000010) && ({row_reg, col_reg}<22'b0001110101100100010011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110101100100010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==22'b0001110101100100010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0001110101100100010101) && ({row_reg, col_reg}<22'b0001110101100100100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100100100010) && ({row_reg, col_reg}<22'b0001110101100100101001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100100101001) && ({row_reg, col_reg}<22'b0001110101100100110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100100110110) && ({row_reg, col_reg}<22'b0001110101100100111101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100100111101) && ({row_reg, col_reg}<22'b0001110101100101001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100101001010) && ({row_reg, col_reg}<22'b0001110101100101010001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100101010001) && ({row_reg, col_reg}<22'b0001110101100101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100101011110) && ({row_reg, col_reg}<22'b0001110101100101100101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100101100101) && ({row_reg, col_reg}<22'b0001110101100101110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100101110010) && ({row_reg, col_reg}<22'b0001110101100101111001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100101111001) && ({row_reg, col_reg}<22'b0001110101100110000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100110000110) && ({row_reg, col_reg}<22'b0001110101100110001101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100110001101) && ({row_reg, col_reg}<22'b0001110101100110011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100110011010) && ({row_reg, col_reg}<22'b0001110101100110100001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100110100001) && ({row_reg, col_reg}<22'b0001110101100110101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100110101110) && ({row_reg, col_reg}<22'b0001110101100110110101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100110110101) && ({row_reg, col_reg}<22'b0001110101100111000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101100111000010) && ({row_reg, col_reg}<22'b0001110101100111001001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100111001001) && ({row_reg, col_reg}<22'b0001110101100111010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b0001110101100111010110)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101100111010111) && ({row_reg, col_reg}<22'b0001110101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101000000010) && ({row_reg, col_reg}<22'b0001110101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110101101010000010) && ({row_reg, col_reg}<22'b0001110101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101101010101100)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=22'b0001110101101010101101) && ({row_reg, col_reg}<22'b0001110101101010110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101010110010) && ({row_reg, col_reg}<22'b0001110101101010111001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101010111001) && ({row_reg, col_reg}<22'b0001110101101011000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101011000110) && ({row_reg, col_reg}<22'b0001110101101011001101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101011001101) && ({row_reg, col_reg}<22'b0001110101101011011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101011011010) && ({row_reg, col_reg}<22'b0001110101101011100001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101011100001) && ({row_reg, col_reg}<22'b0001110101101011101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101011101110) && ({row_reg, col_reg}<22'b0001110101101011110101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101011110101) && ({row_reg, col_reg}<22'b0001110101101100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101100000010) && ({row_reg, col_reg}<22'b0001110101101100001001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101100001001) && ({row_reg, col_reg}<22'b0001110101101100010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101100010110) && ({row_reg, col_reg}<22'b0001110101101100011101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101100011101) && ({row_reg, col_reg}<22'b0001110101101100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101100101010) && ({row_reg, col_reg}<22'b0001110101101100110001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101100110001) && ({row_reg, col_reg}<22'b0001110101101100111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101100111110) && ({row_reg, col_reg}<22'b0001110101101101000101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101101000101) && ({row_reg, col_reg}<22'b0001110101101101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101101010010) && ({row_reg, col_reg}<22'b0001110101101101011001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110101101101011001) && ({row_reg, col_reg}<22'b0001110101101101100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110101101101100110) && ({row_reg, col_reg}<22'b0001110101101101101101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==22'b0001110101101101101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b0001110101101101101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0001110101101101101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0001110101101101110000) && ({row_reg, col_reg}<22'b0001110101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110101110000000010) && ({row_reg, col_reg}<22'b0001110101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110101110000101101) && ({row_reg, col_reg}<22'b0001110110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110110000001010111) && ({row_reg, col_reg}<22'b0001110110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001110110000010000010) && ({row_reg, col_reg}<22'b0001110110000100010000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110110000100010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110110000100010001) && ({row_reg, col_reg}<22'b0001110110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110110001000000010) && ({row_reg, col_reg}<22'b0001110110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110110001010000010) && ({row_reg, col_reg}<22'b0001110110001101110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110001101110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b0001110110001101110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0001110110001101110100) && ({row_reg, col_reg}<22'b0001110110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110110010000000010) && ({row_reg, col_reg}<22'b0001110110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110110010000101101) && ({row_reg, col_reg}<22'b0001110110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110110100001010111) && ({row_reg, col_reg}<22'b0001110110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001110110100010000010) && ({row_reg, col_reg}<22'b0001110110100100001101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110110100100001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==22'b0001110110100100001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0001110110100100001111) && ({row_reg, col_reg}<22'b0001110110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001110110101000000010) && ({row_reg, col_reg}<22'b0001110110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110110101010000010) && ({row_reg, col_reg}<22'b0001110110101101110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110101101110101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=22'b0001110110101101110110) && ({row_reg, col_reg}<22'b0001110110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110110110000000010) && ({row_reg, col_reg}<22'b0001110110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110110110000101101) && ({row_reg, col_reg}<22'b0001110111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110111000001010111) && ({row_reg, col_reg}<22'b0001110111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110111000010000010) && ({row_reg, col_reg}<22'b0001110111000100001100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110111000100001100)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0001110111000100001101) && ({row_reg, col_reg}<22'b0001110111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001110111001000000010) && ({row_reg, col_reg}<22'b0001110111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110111001010000010) && ({row_reg, col_reg}<22'b0001110111001101110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111001101110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0001110111001101111000) && ({row_reg, col_reg}<22'b0001110111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110111010000000010) && ({row_reg, col_reg}<22'b0001110111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110111010000101101) && ({row_reg, col_reg}<22'b0001110111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001110111100001010111) && ({row_reg, col_reg}<22'b0001110111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001110111100010000010) && ({row_reg, col_reg}<22'b0001110111100100001010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110111100100001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110111100100001011) && ({row_reg, col_reg}<22'b0001110111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001110111101000000010) && ({row_reg, col_reg}<22'b0001110111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110111101010000010) && ({row_reg, col_reg}<22'b0001110111101101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111101101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0001110111101101111001) && ({row_reg, col_reg}<22'b0001110111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001110111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001110111110000000010) && ({row_reg, col_reg}<22'b0001110111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001110111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001110111110000101101) && ({row_reg, col_reg}<22'b0001111000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111000000001010111) && ({row_reg, col_reg}<22'b0001111000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001111000000010000010) && ({row_reg, col_reg}<22'b0001111000000100001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111000000100001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0001111000000100001010) && ({row_reg, col_reg}<22'b0001111000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111000001000000010) && ({row_reg, col_reg}<22'b0001111000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111000001010000010) && ({row_reg, col_reg}<22'b0001111000001101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0001111000001101111010) && ({row_reg, col_reg}<22'b0001111000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111000010000000010) && ({row_reg, col_reg}<22'b0001111000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111000010000101101) && ({row_reg, col_reg}<22'b0001111000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111000100001010111) && ({row_reg, col_reg}<22'b0001111000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001111000100010000010) && ({row_reg, col_reg}<22'b0001111000100100001000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111000100100001000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0001111000100100001001) && ({row_reg, col_reg}<22'b0001111000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111000101000000010) && ({row_reg, col_reg}<22'b0001111000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111000101010000010) && ({row_reg, col_reg}<22'b0001111000101101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111000101101111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111000101101111100) && ({row_reg, col_reg}<22'b0001111000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111000110000000010) && ({row_reg, col_reg}<22'b0001111000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111000110000101101) && ({row_reg, col_reg}<22'b0001111001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111001000001010111) && ({row_reg, col_reg}<22'b0001111001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001111001000010000010) && ({row_reg, col_reg}<22'b0001111001000100000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111001000100000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0001111001000100001000) && ({row_reg, col_reg}<22'b0001111001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111001001000000010) && ({row_reg, col_reg}<22'b0001111001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111001001010000010) && ({row_reg, col_reg}<22'b0001111001001101111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0001111001001101111100) && ({row_reg, col_reg}<22'b0001111001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111001010000000010) && ({row_reg, col_reg}<22'b0001111001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111001010000101101) && ({row_reg, col_reg}<22'b0001111001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111001100001010111) && ({row_reg, col_reg}<22'b0001111001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111001100010000010) && ({row_reg, col_reg}<22'b0001111001100100000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111001100100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0001111001100100000111) && ({row_reg, col_reg}<22'b0001111001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111001101000000010) && ({row_reg, col_reg}<22'b0001111001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111001101010000010) && ({row_reg, col_reg}<22'b0001111001101101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0001111001101101111101) && ({row_reg, col_reg}<22'b0001111001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111001110000000010) && ({row_reg, col_reg}<22'b0001111001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111001110000101101) && ({row_reg, col_reg}<22'b0001111010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111010000001010111) && ({row_reg, col_reg}<22'b0001111010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111010000010000010) && ({row_reg, col_reg}<22'b0001111010000100000101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111010000100000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0001111010000100000110) && ({row_reg, col_reg}<22'b0001111010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111010001000000010) && ({row_reg, col_reg}<22'b0001111010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111010001010000010) && ({row_reg, col_reg}<22'b0001111010001101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010001101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0001111010001101111110) && ({row_reg, col_reg}<22'b0001111010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111010010000000010) && ({row_reg, col_reg}<22'b0001111010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111010010000101101) && ({row_reg, col_reg}<22'b0001111010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111010100001010111) && ({row_reg, col_reg}<22'b0001111010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111010100010000010) && ({row_reg, col_reg}<22'b0001111010100100000101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111010100100000101) && ({row_reg, col_reg}<22'b0001111010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111010101000000010) && ({row_reg, col_reg}<22'b0001111010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111010101010000010) && ({row_reg, col_reg}<22'b0001111010101101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010101101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0001111010101101111111) && ({row_reg, col_reg}<22'b0001111010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111010110000000010) && ({row_reg, col_reg}<22'b0001111010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111010110000101101) && ({row_reg, col_reg}<22'b0001111011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111011000001010111) && ({row_reg, col_reg}<22'b0001111011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111011000010000010) && ({row_reg, col_reg}<22'b0001111011000100000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111011000100000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0001111011000100000101) && ({row_reg, col_reg}<22'b0001111011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111011001000000010) && ({row_reg, col_reg}<22'b0001111011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111011001010000010) && ({row_reg, col_reg}<22'b0001111011001101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0001111011001101111111) && ({row_reg, col_reg}<22'b0001111011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111011010000000010) && ({row_reg, col_reg}<22'b0001111011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111011010000101101) && ({row_reg, col_reg}<22'b0001111011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111011100001010111) && ({row_reg, col_reg}<22'b0001111011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111011100010000010) && ({row_reg, col_reg}<22'b0001111011100100000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111011100100000100) && ({row_reg, col_reg}<22'b0001111011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111011101000000010) && ({row_reg, col_reg}<22'b0001111011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111011101010000010) && ({row_reg, col_reg}<22'b0001111011101101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111011101101111111)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=22'b0001111011101110000000) && ({row_reg, col_reg}<22'b0001111011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111011110000000010) && ({row_reg, col_reg}<22'b0001111011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111011110000101101) && ({row_reg, col_reg}<22'b0001111100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111100000001010111) && ({row_reg, col_reg}<22'b0001111100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111100000010000010) && ({row_reg, col_reg}<22'b0001111100000100000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111100000100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0001111100000100000100) && ({row_reg, col_reg}<22'b0001111100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111100001000000010) && ({row_reg, col_reg}<22'b0001111100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111100001010000010) && ({row_reg, col_reg}<22'b0001111100001110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0001111100001110000000) && ({row_reg, col_reg}<22'b0001111100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111100010000000010) && ({row_reg, col_reg}<22'b0001111100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111100010000101101) && ({row_reg, col_reg}<22'b0001111100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111100100001010111) && ({row_reg, col_reg}<22'b0001111100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111100100010000010) && ({row_reg, col_reg}<22'b0001111100100100000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111100100100000011) && ({row_reg, col_reg}<22'b0001111100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111100101000000010) && ({row_reg, col_reg}<22'b0001111100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111100101010000010) && ({row_reg, col_reg}<22'b0001111100101110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111100101110000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0001111100101110000001) && ({row_reg, col_reg}<22'b0001111100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111100110000000010) && ({row_reg, col_reg}<22'b0001111100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111100110000101101) && ({row_reg, col_reg}<22'b0001111101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111101000001010111) && ({row_reg, col_reg}<22'b0001111101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111101000010000010) && ({row_reg, col_reg}<22'b0001111101000100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111101000100000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0001111101000100000011) && ({row_reg, col_reg}<22'b0001111101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111101001000000010) && ({row_reg, col_reg}<22'b0001111101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111101001010000010) && ({row_reg, col_reg}<22'b0001111101001110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111101001110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0001111101001110000001) && ({row_reg, col_reg}<22'b0001111101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111101010000000010) && ({row_reg, col_reg}<22'b0001111101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111101010000101101) && ({row_reg, col_reg}<22'b0001111101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111101100001010111) && ({row_reg, col_reg}<22'b0001111101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111101100010000010) && ({row_reg, col_reg}<22'b0001111101100100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111101100100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0001111101100100000011) && ({row_reg, col_reg}<22'b0001111101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111101101000000010) && ({row_reg, col_reg}<22'b0001111101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111101101010000010) && ({row_reg, col_reg}<22'b0001111101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0001111101101110000001) && ({row_reg, col_reg}<22'b0001111101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111101110000000010) && ({row_reg, col_reg}<22'b0001111101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111101110000101101) && ({row_reg, col_reg}<22'b0001111110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111110000001010111) && ({row_reg, col_reg}<22'b0001111110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111110000010000010) && ({row_reg, col_reg}<22'b0001111110000100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111110000100000010) && ({row_reg, col_reg}<22'b0001111110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111110001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001111110001000000010) && ({row_reg, col_reg}<22'b0001111110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111110001010000010) && ({row_reg, col_reg}<22'b0001111110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0001111110001110000001) && ({row_reg, col_reg}<22'b0001111110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111110010000000010) && ({row_reg, col_reg}<22'b0001111110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111110010000101101) && ({row_reg, col_reg}<22'b0001111110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111110100001010111) && ({row_reg, col_reg}<22'b0001111110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111110100010000010) && ({row_reg, col_reg}<22'b0001111110100100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111110100100000010) && ({row_reg, col_reg}<22'b0001111110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0001111110101000000010) && ({row_reg, col_reg}<22'b0001111110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111110101010000010) && ({row_reg, col_reg}<22'b0001111110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111110101110000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0001111110101110000010) && ({row_reg, col_reg}<22'b0001111110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111110110000000010) && ({row_reg, col_reg}<22'b0001111110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111110110000101101) && ({row_reg, col_reg}<22'b0001111111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111111000001010111) && ({row_reg, col_reg}<22'b0001111111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111111000010000010) && ({row_reg, col_reg}<22'b0001111111000100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111111000100000010) && ({row_reg, col_reg}<22'b0001111111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001111111001000000010) && ({row_reg, col_reg}<22'b0001111111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111111001010000010) && ({row_reg, col_reg}<22'b0001111111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111001110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0001111111001110000010) && ({row_reg, col_reg}<22'b0001111111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111111010000000010) && ({row_reg, col_reg}<22'b0001111111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111111010000101101) && ({row_reg, col_reg}<22'b0001111111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111111100001010111) && ({row_reg, col_reg}<22'b0001111111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111111100010000010) && ({row_reg, col_reg}<22'b0001111111100100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0001111111100100000010) && ({row_reg, col_reg}<22'b0001111111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0001111111101000000010) && ({row_reg, col_reg}<22'b0001111111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111111101010000010) && ({row_reg, col_reg}<22'b0001111111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0001111111101110000010) && ({row_reg, col_reg}<22'b0001111111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0001111111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0001111111110000000010) && ({row_reg, col_reg}<22'b0001111111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0001111111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0001111111110000101101) && ({row_reg, col_reg}<22'b0010000000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000000000001010111) && ({row_reg, col_reg}<22'b0010000000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010000000000010000010) && ({row_reg, col_reg}<22'b0010000000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000000000100000010) && ({row_reg, col_reg}<22'b0010000000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010000000001000000010) && ({row_reg, col_reg}<22'b0010000000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000000001010000010) && ({row_reg, col_reg}<22'b0010000000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000000001110000010) && ({row_reg, col_reg}<22'b0010000000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000000010000000010) && ({row_reg, col_reg}<22'b0010000000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000000010000101101) && ({row_reg, col_reg}<22'b0010000000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000000100001010111) && ({row_reg, col_reg}<22'b0010000000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010000000100010000010) && ({row_reg, col_reg}<22'b0010000000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000000100100000010) && ({row_reg, col_reg}<22'b0010000000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000000101000000010) && ({row_reg, col_reg}<22'b0010000000101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000000101010000010) && ({row_reg, col_reg}<22'b0010000000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000000101110000010) && ({row_reg, col_reg}<22'b0010000000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000000110000000010) && ({row_reg, col_reg}<22'b0010000000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000000110000101101) && ({row_reg, col_reg}<22'b0010000001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000001000001010111) && ({row_reg, col_reg}<22'b0010000001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010000001000010000010) && ({row_reg, col_reg}<22'b0010000001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000001000100000010) && ({row_reg, col_reg}<22'b0010000001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000001001000000010) && ({row_reg, col_reg}<22'b0010000001001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000001001010000010) && ({row_reg, col_reg}<22'b0010000001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000001001110000010) && ({row_reg, col_reg}<22'b0010000001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000001010000000010) && ({row_reg, col_reg}<22'b0010000001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000001010000101101) && ({row_reg, col_reg}<22'b0010000001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000001100001010111) && ({row_reg, col_reg}<22'b0010000001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010000001100010000010) && ({row_reg, col_reg}<22'b0010000001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000001100100000010) && ({row_reg, col_reg}<22'b0010000001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001101000000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0010000001101000000010) && ({row_reg, col_reg}<22'b0010000001101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000001101010000010) && ({row_reg, col_reg}<22'b0010000001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000001101110000010) && ({row_reg, col_reg}<22'b0010000001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000001110000000010) && ({row_reg, col_reg}<22'b0010000001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000001110000101101) && ({row_reg, col_reg}<22'b0010000010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000010000001010111) && ({row_reg, col_reg}<22'b0010000010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010000010000010000010) && ({row_reg, col_reg}<22'b0010000010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000010000100000010) && ({row_reg, col_reg}<22'b0010000010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000010001000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000010001000000010) && ({row_reg, col_reg}<22'b0010000010001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000010001010000010) && ({row_reg, col_reg}<22'b0010000010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000010001110000010) && ({row_reg, col_reg}<22'b0010000010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000010010000000010) && ({row_reg, col_reg}<22'b0010000010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000010010000101101) && ({row_reg, col_reg}<22'b0010000010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000010100001010111) && ({row_reg, col_reg}<22'b0010000010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010000010100010000010) && ({row_reg, col_reg}<22'b0010000010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000010100100000010) && ({row_reg, col_reg}<22'b0010000010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0010000010101000000001) && ({row_reg, col_reg}<22'b0010000010101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000010101010000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0010000010101010000011) && ({row_reg, col_reg}<22'b0010000010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000010101110000010) && ({row_reg, col_reg}<22'b0010000010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000010110000000010) && ({row_reg, col_reg}<22'b0010000010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000010110000101101) && ({row_reg, col_reg}<22'b0010000011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000011000001010111) && ({row_reg, col_reg}<22'b0010000011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010000011000010000010) && ({row_reg, col_reg}<22'b0010000011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000011000100000010) && ({row_reg, col_reg}<22'b0010000011001000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011001000000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0010000011001000000001) && ({row_reg, col_reg}<22'b0010000011001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000011001010000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0010000011001010000011) && ({row_reg, col_reg}<22'b0010000011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000011001110000010) && ({row_reg, col_reg}<22'b0010000011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000011010000000010) && ({row_reg, col_reg}<22'b0010000011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000011010000101101) && ({row_reg, col_reg}<22'b0010000011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000011100001010111) && ({row_reg, col_reg}<22'b0010000011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000011100010000010) && ({row_reg, col_reg}<22'b0010000011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000011100100000010) && ({row_reg, col_reg}<22'b0010000011101000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011101000000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0010000011101000000001) && ({row_reg, col_reg}<22'b0010000011101010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000011101010000011) && ({row_reg, col_reg}<22'b0010000011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000011101110000010) && ({row_reg, col_reg}<22'b0010000011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000011110000000010) && ({row_reg, col_reg}<22'b0010000011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000011110000101101) && ({row_reg, col_reg}<22'b0010000100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000100000001010111) && ({row_reg, col_reg}<22'b0010000100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000100000010000010) && ({row_reg, col_reg}<22'b0010000100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000100000100000010) && ({row_reg, col_reg}<22'b0010000100001000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0010000100001000000000) && ({row_reg, col_reg}<22'b0010000100001010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000100001010000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0010000100001010000100) && ({row_reg, col_reg}<22'b0010000100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000100001110000010) && ({row_reg, col_reg}<22'b0010000100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000100010000000010) && ({row_reg, col_reg}<22'b0010000100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000100010000101101) && ({row_reg, col_reg}<22'b0010000100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000100100001010111) && ({row_reg, col_reg}<22'b0010000100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000100100010000010) && ({row_reg, col_reg}<22'b0010000100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000100100100000010) && ({row_reg, col_reg}<22'b0010000100100111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000100100111111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0010000100101000000000) && ({row_reg, col_reg}<22'b0010000100101010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000100101010000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0010000100101010000100) && ({row_reg, col_reg}<22'b0010000100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000100101110000010) && ({row_reg, col_reg}<22'b0010000100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000100110000000010) && ({row_reg, col_reg}<22'b0010000100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000100110000101101) && ({row_reg, col_reg}<22'b0010000101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000101000001010111) && ({row_reg, col_reg}<22'b0010000101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000101000010000010) && ({row_reg, col_reg}<22'b0010000101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000101000100000010) && ({row_reg, col_reg}<22'b0010000101000111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0010000101000111111111) && ({row_reg, col_reg}<22'b0010000101001010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000101001010000100) && ({row_reg, col_reg}<22'b0010000101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000101001110000010) && ({row_reg, col_reg}<22'b0010000101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000101010000000010) && ({row_reg, col_reg}<22'b0010000101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000101010000101101) && ({row_reg, col_reg}<22'b0010000101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000101100001010111) && ({row_reg, col_reg}<22'b0010000101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000101100010000010) && ({row_reg, col_reg}<22'b0010000101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000101100100000010) && ({row_reg, col_reg}<22'b0010000101100111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000101100111111110)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010000101100111111111) && ({row_reg, col_reg}<22'b0010000101101010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000101101010000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000101101010000101) && ({row_reg, col_reg}<22'b0010000101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000101101110000010) && ({row_reg, col_reg}<22'b0010000101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000101110000000010) && ({row_reg, col_reg}<22'b0010000101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000101110000101101) && ({row_reg, col_reg}<22'b0010000110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000110000001010111) && ({row_reg, col_reg}<22'b0010000110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000110000010000010) && ({row_reg, col_reg}<22'b0010000110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000110000100000010) && ({row_reg, col_reg}<22'b0010000110000111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0010000110000111111110) && ({row_reg, col_reg}<22'b0010000110001010000101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000110001010000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0010000110001010000110) && ({row_reg, col_reg}<22'b0010000110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000110001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010000110001110000010) && ({row_reg, col_reg}<22'b0010000110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000110010000000010) && ({row_reg, col_reg}<22'b0010000110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000110010000101101) && ({row_reg, col_reg}<22'b0010000110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000110100001010111) && ({row_reg, col_reg}<22'b0010000110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000110100010000010) && ({row_reg, col_reg}<22'b0010000110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000110100100000010) && ({row_reg, col_reg}<22'b0010000110100111111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000110100111111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000110100111111110) && ({row_reg, col_reg}<22'b0010000110101010000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000110101010000110) && ({row_reg, col_reg}<22'b0010000110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010000110101110000010) && ({row_reg, col_reg}<22'b0010000110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000110110000000010) && ({row_reg, col_reg}<22'b0010000110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000110110000101101) && ({row_reg, col_reg}<22'b0010000111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000111000001010111) && ({row_reg, col_reg}<22'b0010000111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000111000010000010) && ({row_reg, col_reg}<22'b0010000111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000111000100000010) && ({row_reg, col_reg}<22'b0010000111000111111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111000111111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0010000111000111111101) && ({row_reg, col_reg}<22'b0010000111001010000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000111001010000111) && ({row_reg, col_reg}<22'b0010000111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010000111001110000010) && ({row_reg, col_reg}<22'b0010000111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000111010000000010) && ({row_reg, col_reg}<22'b0010000111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000111010000101101) && ({row_reg, col_reg}<22'b0010000111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010000111100001010111) && ({row_reg, col_reg}<22'b0010000111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000111100010000010) && ({row_reg, col_reg}<22'b0010000111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000111100100000010) && ({row_reg, col_reg}<22'b0010000111100111111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111100111111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010000111100111111100) && ({row_reg, col_reg}<22'b0010000111101010000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000111101010000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000111101010001000) && ({row_reg, col_reg}<22'b0010000111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010000111101110000010) && ({row_reg, col_reg}<22'b0010000111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010000111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010000111110000000010) && ({row_reg, col_reg}<22'b0010000111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010000111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010000111110000101101) && ({row_reg, col_reg}<22'b0010001000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001000000001010111) && ({row_reg, col_reg}<22'b0010001000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001000000010000010) && ({row_reg, col_reg}<22'b0010001000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001000000100000010) && ({row_reg, col_reg}<22'b0010001000000111111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000000111111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001000000111111011) && ({row_reg, col_reg}<22'b0010001000001010001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001000001010001001) && ({row_reg, col_reg}<22'b0010001000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010001000001110000010) && ({row_reg, col_reg}<22'b0010001000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001000010000000010) && ({row_reg, col_reg}<22'b0010001000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001000010000101101) && ({row_reg, col_reg}<22'b0010001000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001000100001010111) && ({row_reg, col_reg}<22'b0010001000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001000100010000010) && ({row_reg, col_reg}<22'b0010001000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001000100100000010) && ({row_reg, col_reg}<22'b0010001000100111111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000100111111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0010001000100111111010) && ({row_reg, col_reg}<22'b0010001000101010001010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001000101010001010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0010001000101010001011) && ({row_reg, col_reg}<22'b0010001000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010001000101110000010) && ({row_reg, col_reg}<22'b0010001000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001000110000000010) && ({row_reg, col_reg}<22'b0010001000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001000110000101101) && ({row_reg, col_reg}<22'b0010001001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001001000001010111) && ({row_reg, col_reg}<22'b0010001001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001001000010000010) && ({row_reg, col_reg}<22'b0010001001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001001000100000010) && ({row_reg, col_reg}<22'b0010001001000111110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001000111110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0010001001000111111000) && ({row_reg, col_reg}<22'b0010001001001010001011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001001001010001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001001001010001100) && ({row_reg, col_reg}<22'b0010001001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010001001001110000010) && ({row_reg, col_reg}<22'b0010001001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001001010000000010) && ({row_reg, col_reg}<22'b0010001001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001001010000101101) && ({row_reg, col_reg}<22'b0010001001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001001100001010111) && ({row_reg, col_reg}<22'b0010001001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001001100010000010) && ({row_reg, col_reg}<22'b0010001001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001001100100000010) && ({row_reg, col_reg}<22'b0010001001100111110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001100111110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==22'b0010001001100111110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0010001001100111110111) && ({row_reg, col_reg}<22'b0010001001101010001101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001001101010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0010001001101010001110) && ({row_reg, col_reg}<22'b0010001001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001001101110000010) && ({row_reg, col_reg}<22'b0010001001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001001110000000010) && ({row_reg, col_reg}<22'b0010001001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001001110000101101) && ({row_reg, col_reg}<22'b0010001010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001010000001010111) && ({row_reg, col_reg}<22'b0010001010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010001010000010000010) && ({row_reg, col_reg}<22'b0010001010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001010000100000010) && ({row_reg, col_reg}<22'b0010001010000111110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010000111110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b0010001010000111110100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001010000111110101) && ({row_reg, col_reg}<22'b0010001010001010001111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001010001010001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001010001010010000) && ({row_reg, col_reg}<22'b0010001010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001010001110000010) && ({row_reg, col_reg}<22'b0010001010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001010010000000010) && ({row_reg, col_reg}<22'b0010001010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001010010000101101) && ({row_reg, col_reg}<22'b0010001010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001010100001010111) && ({row_reg, col_reg}<22'b0010001010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010001010100010000010) && ({row_reg, col_reg}<22'b0010001010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001010100100000010) && ({row_reg, col_reg}<22'b0010001010100111101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010100111101110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==22'b0010001010100111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b0010001010100111110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0010001010100111110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001010100111110010) && ({row_reg, col_reg}<22'b0010001010101010010010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001010101010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0010001010101010010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b0010001010101010010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0010001010101010010101) && ({row_reg, col_reg}<22'b0010001010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001010101110000010) && ({row_reg, col_reg}<22'b0010001010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001010110000000010) && ({row_reg, col_reg}<22'b0010001010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001010110000101101) && ({row_reg, col_reg}<22'b0010001011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001011000001010111) && ({row_reg, col_reg}<22'b0010001011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010001011000010000010) && ({row_reg, col_reg}<22'b0010001011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001011000100000010) && ({row_reg, col_reg}<22'b0010001011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001011000100101101) && ({row_reg, col_reg}<22'b0010001011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001011001101010111) && ({row_reg, col_reg}<22'b0010001011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001011001110000010) && ({row_reg, col_reg}<22'b0010001011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001011010000000010) && ({row_reg, col_reg}<22'b0010001011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001011010000101101) && ({row_reg, col_reg}<22'b0010001011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001011100001010111) && ({row_reg, col_reg}<22'b0010001011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010001011100010000010) && ({row_reg, col_reg}<22'b0010001011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001011100100000010) && ({row_reg, col_reg}<22'b0010001011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001011100100101101) && ({row_reg, col_reg}<22'b0010001011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001011101101010111) && ({row_reg, col_reg}<22'b0010001011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001011101110000010) && ({row_reg, col_reg}<22'b0010001011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001011110000000010) && ({row_reg, col_reg}<22'b0010001011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001011110000101101) && ({row_reg, col_reg}<22'b0010001100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001100000001010111) && ({row_reg, col_reg}<22'b0010001100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010001100000010000010) && ({row_reg, col_reg}<22'b0010001100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001100000100000010) && ({row_reg, col_reg}<22'b0010001100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001100000100101101) && ({row_reg, col_reg}<22'b0010001100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001100001101010111) && ({row_reg, col_reg}<22'b0010001100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001100001110000010) && ({row_reg, col_reg}<22'b0010001100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001100010000000010) && ({row_reg, col_reg}<22'b0010001100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001100010000101101) && ({row_reg, col_reg}<22'b0010001100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001100100001010111) && ({row_reg, col_reg}<22'b0010001100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010001100100010000010) && ({row_reg, col_reg}<22'b0010001100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001100100100000010) && ({row_reg, col_reg}<22'b0010001100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001100100100101101) && ({row_reg, col_reg}<22'b0010001100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001100101101010111) && ({row_reg, col_reg}<22'b0010001100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001100101110000010) && ({row_reg, col_reg}<22'b0010001100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001100110000000010) && ({row_reg, col_reg}<22'b0010001100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001100110000101101) && ({row_reg, col_reg}<22'b0010001101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001101000001010111) && ({row_reg, col_reg}<22'b0010001101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010001101000010000010) && ({row_reg, col_reg}<22'b0010001101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001101000100000010) && ({row_reg, col_reg}<22'b0010001101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001101000100101101) && ({row_reg, col_reg}<22'b0010001101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001101001101010111) && ({row_reg, col_reg}<22'b0010001101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001101001110000010) && ({row_reg, col_reg}<22'b0010001101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001101010000000010) && ({row_reg, col_reg}<22'b0010001101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001101010000101101) && ({row_reg, col_reg}<22'b0010001101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001101100001010111) && ({row_reg, col_reg}<22'b0010001101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001101100010000010) && ({row_reg, col_reg}<22'b0010001101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001101100100000010) && ({row_reg, col_reg}<22'b0010001101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001101100100101101) && ({row_reg, col_reg}<22'b0010001101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001101101101010111) && ({row_reg, col_reg}<22'b0010001101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001101101110000010) && ({row_reg, col_reg}<22'b0010001101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001101110000000010) && ({row_reg, col_reg}<22'b0010001101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001101110000101101) && ({row_reg, col_reg}<22'b0010001110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001110000001010111) && ({row_reg, col_reg}<22'b0010001110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001110000010000010) && ({row_reg, col_reg}<22'b0010001110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001110000100000010) && ({row_reg, col_reg}<22'b0010001110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001110000100101101) && ({row_reg, col_reg}<22'b0010001110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001110001101010111) && ({row_reg, col_reg}<22'b0010001110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001110001110000010) && ({row_reg, col_reg}<22'b0010001110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001110010000000010) && ({row_reg, col_reg}<22'b0010001110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001110010000101101) && ({row_reg, col_reg}<22'b0010001110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001110100001010111) && ({row_reg, col_reg}<22'b0010001110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001110100010000010) && ({row_reg, col_reg}<22'b0010001110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001110100100000010) && ({row_reg, col_reg}<22'b0010001110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001110100100101101) && ({row_reg, col_reg}<22'b0010001110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001110101101010111) && ({row_reg, col_reg}<22'b0010001110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001110101110000010) && ({row_reg, col_reg}<22'b0010001110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001110110000000010) && ({row_reg, col_reg}<22'b0010001110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001110110000101101) && ({row_reg, col_reg}<22'b0010001111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001111000001010111) && ({row_reg, col_reg}<22'b0010001111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001111000010000010) && ({row_reg, col_reg}<22'b0010001111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001111000100000010) && ({row_reg, col_reg}<22'b0010001111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001111000100101101) && ({row_reg, col_reg}<22'b0010001111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001111001101010111) && ({row_reg, col_reg}<22'b0010001111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001111001110000010) && ({row_reg, col_reg}<22'b0010001111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001111010000000010) && ({row_reg, col_reg}<22'b0010001111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001111010000101101) && ({row_reg, col_reg}<22'b0010001111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001111100001010111) && ({row_reg, col_reg}<22'b0010001111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001111100010000010) && ({row_reg, col_reg}<22'b0010001111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001111100100000010) && ({row_reg, col_reg}<22'b0010001111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001111100100101101) && ({row_reg, col_reg}<22'b0010001111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010001111101101010111) && ({row_reg, col_reg}<22'b0010001111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010001111101110000010) && ({row_reg, col_reg}<22'b0010001111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010001111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010001111110000000010) && ({row_reg, col_reg}<22'b0010001111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010001111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010001111110000101101) && ({row_reg, col_reg}<22'b0010010000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010000000001010111) && ({row_reg, col_reg}<22'b0010010000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010000000010000010) && ({row_reg, col_reg}<22'b0010010000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010000000100000010) && ({row_reg, col_reg}<22'b0010010000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010000000100101101) && ({row_reg, col_reg}<22'b0010010000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010000001101010111) && ({row_reg, col_reg}<22'b0010010000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010000001110000010) && ({row_reg, col_reg}<22'b0010010000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010000010000000010) && ({row_reg, col_reg}<22'b0010010000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010000010000101101) && ({row_reg, col_reg}<22'b0010010000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010000100001010111) && ({row_reg, col_reg}<22'b0010010000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010000100010000010) && ({row_reg, col_reg}<22'b0010010000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010000100100000010) && ({row_reg, col_reg}<22'b0010010000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010000100100101101) && ({row_reg, col_reg}<22'b0010010000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010000101101010111) && ({row_reg, col_reg}<22'b0010010000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010000101110000010) && ({row_reg, col_reg}<22'b0010010000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010000110000000010) && ({row_reg, col_reg}<22'b0010010000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010000110000101101) && ({row_reg, col_reg}<22'b0010010001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010001000001010111) && ({row_reg, col_reg}<22'b0010010001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010001000010000010) && ({row_reg, col_reg}<22'b0010010001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010001000100000010) && ({row_reg, col_reg}<22'b0010010001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010001000100101101) && ({row_reg, col_reg}<22'b0010010001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010001001101010111) && ({row_reg, col_reg}<22'b0010010001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010010001001110000010) && ({row_reg, col_reg}<22'b0010010001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010001010000000010) && ({row_reg, col_reg}<22'b0010010001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010001010000101101) && ({row_reg, col_reg}<22'b0010010001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010001100001010111) && ({row_reg, col_reg}<22'b0010010001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010001100010000010) && ({row_reg, col_reg}<22'b0010010001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010001100100000010) && ({row_reg, col_reg}<22'b0010010001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010001100100101101) && ({row_reg, col_reg}<22'b0010010001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010001101101010111) && ({row_reg, col_reg}<22'b0010010001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010010001101110000010) && ({row_reg, col_reg}<22'b0010010001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010001110000000010) && ({row_reg, col_reg}<22'b0010010001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010001110000101101) && ({row_reg, col_reg}<22'b0010010010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010010000001010111) && ({row_reg, col_reg}<22'b0010010010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010010000010000010) && ({row_reg, col_reg}<22'b0010010010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010010000100000010) && ({row_reg, col_reg}<22'b0010010010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010010000100101101) && ({row_reg, col_reg}<22'b0010010010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010010001101010111) && ({row_reg, col_reg}<22'b0010010010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010010010001110000010) && ({row_reg, col_reg}<22'b0010010010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010010010000000010) && ({row_reg, col_reg}<22'b0010010010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010010010000101101) && ({row_reg, col_reg}<22'b0010010010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010010100001010111) && ({row_reg, col_reg}<22'b0010010010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010010100010000010) && ({row_reg, col_reg}<22'b0010010010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010010100100000010) && ({row_reg, col_reg}<22'b0010010010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010010100100101101) && ({row_reg, col_reg}<22'b0010010010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010010101101010111) && ({row_reg, col_reg}<22'b0010010010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010010101110000010) && ({row_reg, col_reg}<22'b0010010010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010010110000000010) && ({row_reg, col_reg}<22'b0010010010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010010110000101101) && ({row_reg, col_reg}<22'b0010010011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010011000001010111) && ({row_reg, col_reg}<22'b0010010011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010011000010000010) && ({row_reg, col_reg}<22'b0010010011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010011000100000010) && ({row_reg, col_reg}<22'b0010010011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010011000100101101) && ({row_reg, col_reg}<22'b0010010011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010011001101010111) && ({row_reg, col_reg}<22'b0010010011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010011001110000010) && ({row_reg, col_reg}<22'b0010010011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010011010000000010) && ({row_reg, col_reg}<22'b0010010011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010011010000101101) && ({row_reg, col_reg}<22'b0010010011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010011100001010111) && ({row_reg, col_reg}<22'b0010010011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010011100010000010) && ({row_reg, col_reg}<22'b0010010011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010011100100000010) && ({row_reg, col_reg}<22'b0010010011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010011100100101101) && ({row_reg, col_reg}<22'b0010010011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010011101101010111) && ({row_reg, col_reg}<22'b0010010011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010011101110000010) && ({row_reg, col_reg}<22'b0010010011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010011110000000010) && ({row_reg, col_reg}<22'b0010010011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010011110000101101) && ({row_reg, col_reg}<22'b0010010100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010100000001010111) && ({row_reg, col_reg}<22'b0010010100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010100000010000010) && ({row_reg, col_reg}<22'b0010010100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010100000100000010) && ({row_reg, col_reg}<22'b0010010100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010100000100101101) && ({row_reg, col_reg}<22'b0010010100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010100001101010111) && ({row_reg, col_reg}<22'b0010010100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010100001110000010) && ({row_reg, col_reg}<22'b0010010100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010100010000000010) && ({row_reg, col_reg}<22'b0010010100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010100010000101101) && ({row_reg, col_reg}<22'b0010010100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010100100001010111) && ({row_reg, col_reg}<22'b0010010100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010100100010000010) && ({row_reg, col_reg}<22'b0010010100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010100100100000010) && ({row_reg, col_reg}<22'b0010010100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010100100100101101) && ({row_reg, col_reg}<22'b0010010100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010100101101010111) && ({row_reg, col_reg}<22'b0010010100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010100101110000010) && ({row_reg, col_reg}<22'b0010010100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010100110000000010) && ({row_reg, col_reg}<22'b0010010100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010100110000101101) && ({row_reg, col_reg}<22'b0010010101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010101000001010111) && ({row_reg, col_reg}<22'b0010010101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010010101000010000010) && ({row_reg, col_reg}<22'b0010010101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010101000100000010) && ({row_reg, col_reg}<22'b0010010101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010101000100101101) && ({row_reg, col_reg}<22'b0010010101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010101001101010111) && ({row_reg, col_reg}<22'b0010010101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010101001110000010) && ({row_reg, col_reg}<22'b0010010101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010101010000000010) && ({row_reg, col_reg}<22'b0010010101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010101010000101101) && ({row_reg, col_reg}<22'b0010010101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010101100001010111) && ({row_reg, col_reg}<22'b0010010101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010010101100010000010) && ({row_reg, col_reg}<22'b0010010101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010101100100000010) && ({row_reg, col_reg}<22'b0010010101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010101100100101101) && ({row_reg, col_reg}<22'b0010010101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010101101101010111) && ({row_reg, col_reg}<22'b0010010101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010101101110000010) && ({row_reg, col_reg}<22'b0010010101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010101110000000010) && ({row_reg, col_reg}<22'b0010010101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010101110000101101) && ({row_reg, col_reg}<22'b0010010110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010110000001010111) && ({row_reg, col_reg}<22'b0010010110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010010110000010000010) && ({row_reg, col_reg}<22'b0010010110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010110000100000010) && ({row_reg, col_reg}<22'b0010010110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010110000100101101) && ({row_reg, col_reg}<22'b0010010110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010110001101010111) && ({row_reg, col_reg}<22'b0010010110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010110001110000010) && ({row_reg, col_reg}<22'b0010010110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010110010000000010) && ({row_reg, col_reg}<22'b0010010110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010110010000101101) && ({row_reg, col_reg}<22'b0010010110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010110100001010111) && ({row_reg, col_reg}<22'b0010010110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010110100010000010) && ({row_reg, col_reg}<22'b0010010110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010110100100000010) && ({row_reg, col_reg}<22'b0010010110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010110100100101101) && ({row_reg, col_reg}<22'b0010010110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010110101101010111) && ({row_reg, col_reg}<22'b0010010110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010110101110000010) && ({row_reg, col_reg}<22'b0010010110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010110110000000010) && ({row_reg, col_reg}<22'b0010010110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010110110000101101) && ({row_reg, col_reg}<22'b0010010111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010111000001010111) && ({row_reg, col_reg}<22'b0010010111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010010111000010000010) && ({row_reg, col_reg}<22'b0010010111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010111000100000010) && ({row_reg, col_reg}<22'b0010010111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010111000100101101) && ({row_reg, col_reg}<22'b0010010111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010111001101010111) && ({row_reg, col_reg}<22'b0010010111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010111001110000010) && ({row_reg, col_reg}<22'b0010010111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010111010000000010) && ({row_reg, col_reg}<22'b0010010111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010111010000101101) && ({row_reg, col_reg}<22'b0010010111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010111100001010111) && ({row_reg, col_reg}<22'b0010010111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010111100010000010) && ({row_reg, col_reg}<22'b0010010111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010111100100000010) && ({row_reg, col_reg}<22'b0010010111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010111100100101101) && ({row_reg, col_reg}<22'b0010010111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010010111101101010111) && ({row_reg, col_reg}<22'b0010010111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010010111101110000010) && ({row_reg, col_reg}<22'b0010010111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010010111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010010111110000000010) && ({row_reg, col_reg}<22'b0010010111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010010111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010010111110000101101) && ({row_reg, col_reg}<22'b0010011000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011000000001010111) && ({row_reg, col_reg}<22'b0010011000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011000000010000010) && ({row_reg, col_reg}<22'b0010011000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011000000100000010) && ({row_reg, col_reg}<22'b0010011000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011000000100101101) && ({row_reg, col_reg}<22'b0010011000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011000001101010111) && ({row_reg, col_reg}<22'b0010011000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011000001110000010) && ({row_reg, col_reg}<22'b0010011000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011000010000000010) && ({row_reg, col_reg}<22'b0010011000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011000010000101101) && ({row_reg, col_reg}<22'b0010011000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011000100001010111) && ({row_reg, col_reg}<22'b0010011000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011000100010000010) && ({row_reg, col_reg}<22'b0010011000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011000100100000010) && ({row_reg, col_reg}<22'b0010011000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011000100100101101) && ({row_reg, col_reg}<22'b0010011000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011000101101010111) && ({row_reg, col_reg}<22'b0010011000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011000101110000010) && ({row_reg, col_reg}<22'b0010011000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011000110000000010) && ({row_reg, col_reg}<22'b0010011000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011000110000101101) && ({row_reg, col_reg}<22'b0010011001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011001000001010111) && ({row_reg, col_reg}<22'b0010011001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011001000010000010) && ({row_reg, col_reg}<22'b0010011001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011001000100000010) && ({row_reg, col_reg}<22'b0010011001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011001000100101101) && ({row_reg, col_reg}<22'b0010011001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011001001101010111) && ({row_reg, col_reg}<22'b0010011001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011001001110000010) && ({row_reg, col_reg}<22'b0010011001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011001010000000010) && ({row_reg, col_reg}<22'b0010011001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011001010000101101) && ({row_reg, col_reg}<22'b0010011001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011001100001010111) && ({row_reg, col_reg}<22'b0010011001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011001100010000010) && ({row_reg, col_reg}<22'b0010011001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011001100100000010) && ({row_reg, col_reg}<22'b0010011001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011001100100101101) && ({row_reg, col_reg}<22'b0010011001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011001101101010111) && ({row_reg, col_reg}<22'b0010011001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011001101110000010) && ({row_reg, col_reg}<22'b0010011001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011001110000000010) && ({row_reg, col_reg}<22'b0010011001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011001110000101101) && ({row_reg, col_reg}<22'b0010011010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011010000001010111) && ({row_reg, col_reg}<22'b0010011010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011010000010000010) && ({row_reg, col_reg}<22'b0010011010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011010000100000010) && ({row_reg, col_reg}<22'b0010011010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011010000100101101) && ({row_reg, col_reg}<22'b0010011010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011010001101010111) && ({row_reg, col_reg}<22'b0010011010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010011010001110000010) && ({row_reg, col_reg}<22'b0010011010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011010010000000010) && ({row_reg, col_reg}<22'b0010011010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011010010000101101) && ({row_reg, col_reg}<22'b0010011010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011010100001010111) && ({row_reg, col_reg}<22'b0010011010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011010100010000010) && ({row_reg, col_reg}<22'b0010011010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011010100100000010) && ({row_reg, col_reg}<22'b0010011010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011010100100101101) && ({row_reg, col_reg}<22'b0010011010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011010101101010111) && ({row_reg, col_reg}<22'b0010011010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010011010101110000010) && ({row_reg, col_reg}<22'b0010011010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011010110000000010) && ({row_reg, col_reg}<22'b0010011010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011010110000101101) && ({row_reg, col_reg}<22'b0010011011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011011000001010111) && ({row_reg, col_reg}<22'b0010011011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011011000010000010) && ({row_reg, col_reg}<22'b0010011011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011011000100000010) && ({row_reg, col_reg}<22'b0010011011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011011000100101101) && ({row_reg, col_reg}<22'b0010011011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011011001101010111) && ({row_reg, col_reg}<22'b0010011011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010011011001110000010) && ({row_reg, col_reg}<22'b0010011011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011011010000000010) && ({row_reg, col_reg}<22'b0010011011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011011010000101101) && ({row_reg, col_reg}<22'b0010011011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011011100001010111) && ({row_reg, col_reg}<22'b0010011011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011011100010000010) && ({row_reg, col_reg}<22'b0010011011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011011100100000010) && ({row_reg, col_reg}<22'b0010011011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011011100100101101) && ({row_reg, col_reg}<22'b0010011011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011011101101010111) && ({row_reg, col_reg}<22'b0010011011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010011011101110000010) && ({row_reg, col_reg}<22'b0010011011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011011110000000010) && ({row_reg, col_reg}<22'b0010011011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011011110000101101) && ({row_reg, col_reg}<22'b0010011100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011100000001010111) && ({row_reg, col_reg}<22'b0010011100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011100000010000010) && ({row_reg, col_reg}<22'b0010011100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011100000100000010) && ({row_reg, col_reg}<22'b0010011100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011100000100101101) && ({row_reg, col_reg}<22'b0010011100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011100001101010111) && ({row_reg, col_reg}<22'b0010011100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010011100001110000010) && ({row_reg, col_reg}<22'b0010011100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011100010000000010) && ({row_reg, col_reg}<22'b0010011100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011100010000101101) && ({row_reg, col_reg}<22'b0010011100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011100100001010111) && ({row_reg, col_reg}<22'b0010011100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011100100010000010) && ({row_reg, col_reg}<22'b0010011100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011100100100000010) && ({row_reg, col_reg}<22'b0010011100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011100100100101101) && ({row_reg, col_reg}<22'b0010011100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011100101101010111) && ({row_reg, col_reg}<22'b0010011100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010011100101110000010) && ({row_reg, col_reg}<22'b0010011100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011100110000000010) && ({row_reg, col_reg}<22'b0010011100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011100110000101101) && ({row_reg, col_reg}<22'b0010011101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011101000001010111) && ({row_reg, col_reg}<22'b0010011101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011101000010000010) && ({row_reg, col_reg}<22'b0010011101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011101000100000010) && ({row_reg, col_reg}<22'b0010011101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011101000100101101) && ({row_reg, col_reg}<22'b0010011101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011101001101010111) && ({row_reg, col_reg}<22'b0010011101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010011101001110000010) && ({row_reg, col_reg}<22'b0010011101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011101010000000010) && ({row_reg, col_reg}<22'b0010011101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011101010000101101) && ({row_reg, col_reg}<22'b0010011101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011101100001010111) && ({row_reg, col_reg}<22'b0010011101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011101100010000010) && ({row_reg, col_reg}<22'b0010011101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011101100100000010) && ({row_reg, col_reg}<22'b0010011101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011101100100101101) && ({row_reg, col_reg}<22'b0010011101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011101101101010111) && ({row_reg, col_reg}<22'b0010011101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011101101110000010) && ({row_reg, col_reg}<22'b0010011101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011101110000000010) && ({row_reg, col_reg}<22'b0010011101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011101110000101101) && ({row_reg, col_reg}<22'b0010011110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011110000001010111) && ({row_reg, col_reg}<22'b0010011110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010011110000010000010) && ({row_reg, col_reg}<22'b0010011110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011110000100000010) && ({row_reg, col_reg}<22'b0010011110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011110000100101101) && ({row_reg, col_reg}<22'b0010011110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011110001101010111) && ({row_reg, col_reg}<22'b0010011110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011110001110000010) && ({row_reg, col_reg}<22'b0010011110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011110010000000010) && ({row_reg, col_reg}<22'b0010011110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011110010000101101) && ({row_reg, col_reg}<22'b0010011110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011110100001010111) && ({row_reg, col_reg}<22'b0010011110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010011110100010000010) && ({row_reg, col_reg}<22'b0010011110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011110100100000010) && ({row_reg, col_reg}<22'b0010011110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011110100100101101) && ({row_reg, col_reg}<22'b0010011110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011110101101010111) && ({row_reg, col_reg}<22'b0010011110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011110101110000010) && ({row_reg, col_reg}<22'b0010011110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011110110000000010) && ({row_reg, col_reg}<22'b0010011110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011110110000101101) && ({row_reg, col_reg}<22'b0010011111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011111000001010111) && ({row_reg, col_reg}<22'b0010011111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010011111000010000010) && ({row_reg, col_reg}<22'b0010011111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011111000100000010) && ({row_reg, col_reg}<22'b0010011111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011111000100101101) && ({row_reg, col_reg}<22'b0010011111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011111001101010111) && ({row_reg, col_reg}<22'b0010011111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011111001110000010) && ({row_reg, col_reg}<22'b0010011111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011111010000000010) && ({row_reg, col_reg}<22'b0010011111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011111010000101101) && ({row_reg, col_reg}<22'b0010011111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011111100001010111) && ({row_reg, col_reg}<22'b0010011111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010011111100010000010) && ({row_reg, col_reg}<22'b0010011111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011111100100000010) && ({row_reg, col_reg}<22'b0010011111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011111100100101101) && ({row_reg, col_reg}<22'b0010011111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010011111101101010111) && ({row_reg, col_reg}<22'b0010011111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010011111101110000010) && ({row_reg, col_reg}<22'b0010011111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010011111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010011111110000000010) && ({row_reg, col_reg}<22'b0010011111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010011111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010011111110000101101) && ({row_reg, col_reg}<22'b0010100000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100000000001010111) && ({row_reg, col_reg}<22'b0010100000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010100000000010000010) && ({row_reg, col_reg}<22'b0010100000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100000000100000010) && ({row_reg, col_reg}<22'b0010100000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100000000100101101) && ({row_reg, col_reg}<22'b0010100000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100000001101010111) && ({row_reg, col_reg}<22'b0010100000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100000001110000010) && ({row_reg, col_reg}<22'b0010100000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100000010000000010) && ({row_reg, col_reg}<22'b0010100000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100000010000101101) && ({row_reg, col_reg}<22'b0010100000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100000100001010111) && ({row_reg, col_reg}<22'b0010100000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010100000100010000010) && ({row_reg, col_reg}<22'b0010100000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100000100100000010) && ({row_reg, col_reg}<22'b0010100000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100000100100101101) && ({row_reg, col_reg}<22'b0010100000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100000101101010111) && ({row_reg, col_reg}<22'b0010100000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100000101110000010) && ({row_reg, col_reg}<22'b0010100000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100000110000000010) && ({row_reg, col_reg}<22'b0010100000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100000110000101101) && ({row_reg, col_reg}<22'b0010100001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100001000001010111) && ({row_reg, col_reg}<22'b0010100001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010100001000010000010) && ({row_reg, col_reg}<22'b0010100001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100001000100000010) && ({row_reg, col_reg}<22'b0010100001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100001000100101101) && ({row_reg, col_reg}<22'b0010100001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100001001101010111) && ({row_reg, col_reg}<22'b0010100001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100001001110000010) && ({row_reg, col_reg}<22'b0010100001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100001010000000010) && ({row_reg, col_reg}<22'b0010100001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100001010000101101) && ({row_reg, col_reg}<22'b0010100001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100001100001010111) && ({row_reg, col_reg}<22'b0010100001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100001100010000010) && ({row_reg, col_reg}<22'b0010100001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100001100100000010) && ({row_reg, col_reg}<22'b0010100001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100001100100101101) && ({row_reg, col_reg}<22'b0010100001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100001101101010111) && ({row_reg, col_reg}<22'b0010100001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100001101110000010) && ({row_reg, col_reg}<22'b0010100001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100001110000000010) && ({row_reg, col_reg}<22'b0010100001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100001110000101101) && ({row_reg, col_reg}<22'b0010100010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100010000001010111) && ({row_reg, col_reg}<22'b0010100010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100010000010000010) && ({row_reg, col_reg}<22'b0010100010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100010000100000010) && ({row_reg, col_reg}<22'b0010100010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100010000100101101) && ({row_reg, col_reg}<22'b0010100010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100010001101010111) && ({row_reg, col_reg}<22'b0010100010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100010001110000010) && ({row_reg, col_reg}<22'b0010100010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100010010000000010) && ({row_reg, col_reg}<22'b0010100010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100010010000101101) && ({row_reg, col_reg}<22'b0010100010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100010100001010111) && ({row_reg, col_reg}<22'b0010100010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100010100010000010) && ({row_reg, col_reg}<22'b0010100010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100010100100000010) && ({row_reg, col_reg}<22'b0010100010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100010100100101101) && ({row_reg, col_reg}<22'b0010100010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100010101101010111) && ({row_reg, col_reg}<22'b0010100010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100010101110000010) && ({row_reg, col_reg}<22'b0010100010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100010110000000010) && ({row_reg, col_reg}<22'b0010100010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100010110000101101) && ({row_reg, col_reg}<22'b0010100011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100011000001010111) && ({row_reg, col_reg}<22'b0010100011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100011000010000010) && ({row_reg, col_reg}<22'b0010100011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100011000100000010) && ({row_reg, col_reg}<22'b0010100011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100011000100101101) && ({row_reg, col_reg}<22'b0010100011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100011001101010111) && ({row_reg, col_reg}<22'b0010100011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100011001110000010) && ({row_reg, col_reg}<22'b0010100011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100011010000000010) && ({row_reg, col_reg}<22'b0010100011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100011010000101101) && ({row_reg, col_reg}<22'b0010100011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100011100001010111) && ({row_reg, col_reg}<22'b0010100011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100011100010000010) && ({row_reg, col_reg}<22'b0010100011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100011100100000010) && ({row_reg, col_reg}<22'b0010100011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100011100100101101) && ({row_reg, col_reg}<22'b0010100011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100011101101010111) && ({row_reg, col_reg}<22'b0010100011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100011101110000010) && ({row_reg, col_reg}<22'b0010100011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100011110000000010) && ({row_reg, col_reg}<22'b0010100011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100011110000101101) && ({row_reg, col_reg}<22'b0010100100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100100000001010111) && ({row_reg, col_reg}<22'b0010100100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100100000010000010) && ({row_reg, col_reg}<22'b0010100100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100100000100000010) && ({row_reg, col_reg}<22'b0010100100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100100000100101101) && ({row_reg, col_reg}<22'b0010100100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100100001101010111) && ({row_reg, col_reg}<22'b0010100100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010100100001110000010) && ({row_reg, col_reg}<22'b0010100100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100100010000000010) && ({row_reg, col_reg}<22'b0010100100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100100010000101101) && ({row_reg, col_reg}<22'b0010100100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100100100001010111) && ({row_reg, col_reg}<22'b0010100100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100100100010000010) && ({row_reg, col_reg}<22'b0010100100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100100100100000010) && ({row_reg, col_reg}<22'b0010100100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100100100100101101) && ({row_reg, col_reg}<22'b0010100100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100100101101010111) && ({row_reg, col_reg}<22'b0010100100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010100100101110000010) && ({row_reg, col_reg}<22'b0010100100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100100110000000010) && ({row_reg, col_reg}<22'b0010100100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100100110000101101) && ({row_reg, col_reg}<22'b0010100101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100101000001010111) && ({row_reg, col_reg}<22'b0010100101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100101000010000010) && ({row_reg, col_reg}<22'b0010100101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100101000100000010) && ({row_reg, col_reg}<22'b0010100101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100101000100101101) && ({row_reg, col_reg}<22'b0010100101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100101001101010111) && ({row_reg, col_reg}<22'b0010100101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010100101001110000010) && ({row_reg, col_reg}<22'b0010100101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100101010000000010) && ({row_reg, col_reg}<22'b0010100101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100101010000101101) && ({row_reg, col_reg}<22'b0010100101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100101100001010111) && ({row_reg, col_reg}<22'b0010100101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100101100010000010) && ({row_reg, col_reg}<22'b0010100101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100101100100000010) && ({row_reg, col_reg}<22'b0010100101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100101100100101101) && ({row_reg, col_reg}<22'b0010100101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100101101101010111) && ({row_reg, col_reg}<22'b0010100101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010100101101110000010) && ({row_reg, col_reg}<22'b0010100101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100101110000000010) && ({row_reg, col_reg}<22'b0010100101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100101110000101101) && ({row_reg, col_reg}<22'b0010100110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100110000001010111) && ({row_reg, col_reg}<22'b0010100110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100110000010000010) && ({row_reg, col_reg}<22'b0010100110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100110000100000010) && ({row_reg, col_reg}<22'b0010100110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100110000100101101) && ({row_reg, col_reg}<22'b0010100110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100110001101010111) && ({row_reg, col_reg}<22'b0010100110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010100110001110000010) && ({row_reg, col_reg}<22'b0010100110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100110010000000010) && ({row_reg, col_reg}<22'b0010100110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100110010000101101) && ({row_reg, col_reg}<22'b0010100110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100110100001010111) && ({row_reg, col_reg}<22'b0010100110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100110100010000010) && ({row_reg, col_reg}<22'b0010100110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100110100100000010) && ({row_reg, col_reg}<22'b0010100110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100110100100101101) && ({row_reg, col_reg}<22'b0010100110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100110101101010111) && ({row_reg, col_reg}<22'b0010100110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010100110101110000010) && ({row_reg, col_reg}<22'b0010100110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100110110000000010) && ({row_reg, col_reg}<22'b0010100110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100110110000101101) && ({row_reg, col_reg}<22'b0010100111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100111000001010111) && ({row_reg, col_reg}<22'b0010100111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100111000010000010) && ({row_reg, col_reg}<22'b0010100111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100111000100000010) && ({row_reg, col_reg}<22'b0010100111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100111000100101101) && ({row_reg, col_reg}<22'b0010100111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100111001101010111) && ({row_reg, col_reg}<22'b0010100111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010100111001110000010) && ({row_reg, col_reg}<22'b0010100111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100111010000000010) && ({row_reg, col_reg}<22'b0010100111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100111010000101101) && ({row_reg, col_reg}<22'b0010100111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100111100001010111) && ({row_reg, col_reg}<22'b0010100111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100111100010000010) && ({row_reg, col_reg}<22'b0010100111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100111100100000010) && ({row_reg, col_reg}<22'b0010100111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100111100100101101) && ({row_reg, col_reg}<22'b0010100111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010100111101101010111) && ({row_reg, col_reg}<22'b0010100111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010100111101110000010) && ({row_reg, col_reg}<22'b0010100111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010100111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010100111110000000010) && ({row_reg, col_reg}<22'b0010100111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010100111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010100111110000101101) && ({row_reg, col_reg}<22'b0010101000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101000000001010111) && ({row_reg, col_reg}<22'b0010101000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010101000000010000010) && ({row_reg, col_reg}<22'b0010101000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101000000100000010) && ({row_reg, col_reg}<22'b0010101000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101000000100101101) && ({row_reg, col_reg}<22'b0010101000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101000001101010111) && ({row_reg, col_reg}<22'b0010101000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101000001110000010) && ({row_reg, col_reg}<22'b0010101000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101000010000000010) && ({row_reg, col_reg}<22'b0010101000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101000010000101101) && ({row_reg, col_reg}<22'b0010101000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101000100001010111) && ({row_reg, col_reg}<22'b0010101000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010101000100010000010) && ({row_reg, col_reg}<22'b0010101000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101000100100000010) && ({row_reg, col_reg}<22'b0010101000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101000100100101101) && ({row_reg, col_reg}<22'b0010101000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101000101101010111) && ({row_reg, col_reg}<22'b0010101000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101000101110000010) && ({row_reg, col_reg}<22'b0010101000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101000110000000010) && ({row_reg, col_reg}<22'b0010101000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101000110000101101) && ({row_reg, col_reg}<22'b0010101001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101001000001010111) && ({row_reg, col_reg}<22'b0010101001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010101001000010000010) && ({row_reg, col_reg}<22'b0010101001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101001000100000010) && ({row_reg, col_reg}<22'b0010101001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101001000100101101) && ({row_reg, col_reg}<22'b0010101001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101001001101010111) && ({row_reg, col_reg}<22'b0010101001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101001001110000010) && ({row_reg, col_reg}<22'b0010101001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101001010000000010) && ({row_reg, col_reg}<22'b0010101001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101001010000101101) && ({row_reg, col_reg}<22'b0010101001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101001100001010111) && ({row_reg, col_reg}<22'b0010101001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010101001100010000010) && ({row_reg, col_reg}<22'b0010101001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101001100100000010) && ({row_reg, col_reg}<22'b0010101001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101001100100101101) && ({row_reg, col_reg}<22'b0010101001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101001101101010111) && ({row_reg, col_reg}<22'b0010101001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101001101110000010) && ({row_reg, col_reg}<22'b0010101001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101001110000000010) && ({row_reg, col_reg}<22'b0010101001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101001110000101101) && ({row_reg, col_reg}<22'b0010101010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101010000001010111) && ({row_reg, col_reg}<22'b0010101010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010101010000010000010) && ({row_reg, col_reg}<22'b0010101010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101010000100000010) && ({row_reg, col_reg}<22'b0010101010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101010000100101101) && ({row_reg, col_reg}<22'b0010101010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101010001101010111) && ({row_reg, col_reg}<22'b0010101010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101010001110000010) && ({row_reg, col_reg}<22'b0010101010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101010010000000010) && ({row_reg, col_reg}<22'b0010101010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101010010000101101) && ({row_reg, col_reg}<22'b0010101010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101010100001010111) && ({row_reg, col_reg}<22'b0010101010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010101010100010000010) && ({row_reg, col_reg}<22'b0010101010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101010100100000010) && ({row_reg, col_reg}<22'b0010101010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101010100100101101) && ({row_reg, col_reg}<22'b0010101010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101010101101010111) && ({row_reg, col_reg}<22'b0010101010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101010101110000010) && ({row_reg, col_reg}<22'b0010101010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101010110000000010) && ({row_reg, col_reg}<22'b0010101010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101010110000101101) && ({row_reg, col_reg}<22'b0010101011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101011000001010111) && ({row_reg, col_reg}<22'b0010101011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010101011000010000010) && ({row_reg, col_reg}<22'b0010101011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101011000100000010) && ({row_reg, col_reg}<22'b0010101011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101011000100101101) && ({row_reg, col_reg}<22'b0010101011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101011001101010111) && ({row_reg, col_reg}<22'b0010101011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101011001110000010) && ({row_reg, col_reg}<22'b0010101011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101011010000000010) && ({row_reg, col_reg}<22'b0010101011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101011010000101101) && ({row_reg, col_reg}<22'b0010101011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101011100001010111) && ({row_reg, col_reg}<22'b0010101011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101011100010000010) && ({row_reg, col_reg}<22'b0010101011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101011100100000010) && ({row_reg, col_reg}<22'b0010101011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101011100100101101) && ({row_reg, col_reg}<22'b0010101011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101011101101010111) && ({row_reg, col_reg}<22'b0010101011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101011101110000010) && ({row_reg, col_reg}<22'b0010101011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101011110000000010) && ({row_reg, col_reg}<22'b0010101011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101011110000101101) && ({row_reg, col_reg}<22'b0010101100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101100000001010111) && ({row_reg, col_reg}<22'b0010101100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101100000010000010) && ({row_reg, col_reg}<22'b0010101100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101100000100000010) && ({row_reg, col_reg}<22'b0010101100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101100000100101101) && ({row_reg, col_reg}<22'b0010101100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101100001101010111) && ({row_reg, col_reg}<22'b0010101100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101100001110000010) && ({row_reg, col_reg}<22'b0010101100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101100010000000010) && ({row_reg, col_reg}<22'b0010101100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101100010000101101) && ({row_reg, col_reg}<22'b0010101100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101100100001010111) && ({row_reg, col_reg}<22'b0010101100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101100100010000010) && ({row_reg, col_reg}<22'b0010101100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101100100100000010) && ({row_reg, col_reg}<22'b0010101100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101100100100101101) && ({row_reg, col_reg}<22'b0010101100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101100101101010111) && ({row_reg, col_reg}<22'b0010101100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101100101110000010) && ({row_reg, col_reg}<22'b0010101100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101100110000000010) && ({row_reg, col_reg}<22'b0010101100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101100110000101101) && ({row_reg, col_reg}<22'b0010101101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101101000001010111) && ({row_reg, col_reg}<22'b0010101101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101101000010000010) && ({row_reg, col_reg}<22'b0010101101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101101000100000010) && ({row_reg, col_reg}<22'b0010101101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101101000100101101) && ({row_reg, col_reg}<22'b0010101101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101101001101010111) && ({row_reg, col_reg}<22'b0010101101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101101001110000010) && ({row_reg, col_reg}<22'b0010101101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101101010000000010) && ({row_reg, col_reg}<22'b0010101101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101101010000101101) && ({row_reg, col_reg}<22'b0010101101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101101100001010111) && ({row_reg, col_reg}<22'b0010101101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101101100010000010) && ({row_reg, col_reg}<22'b0010101101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101101100100000010) && ({row_reg, col_reg}<22'b0010101101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101101100100101101) && ({row_reg, col_reg}<22'b0010101101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101101101101010111) && ({row_reg, col_reg}<22'b0010101101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101101101110000010) && ({row_reg, col_reg}<22'b0010101101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101101110000000010) && ({row_reg, col_reg}<22'b0010101101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101101110000101101) && ({row_reg, col_reg}<22'b0010101110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101110000001010111) && ({row_reg, col_reg}<22'b0010101110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101110000010000010) && ({row_reg, col_reg}<22'b0010101110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101110000100000010) && ({row_reg, col_reg}<22'b0010101110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101110000100101101) && ({row_reg, col_reg}<22'b0010101110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101110001101010111) && ({row_reg, col_reg}<22'b0010101110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010101110001110000010) && ({row_reg, col_reg}<22'b0010101110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101110010000000010) && ({row_reg, col_reg}<22'b0010101110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101110010000101101) && ({row_reg, col_reg}<22'b0010101110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101110100001010111) && ({row_reg, col_reg}<22'b0010101110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101110100010000010) && ({row_reg, col_reg}<22'b0010101110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101110100100000010) && ({row_reg, col_reg}<22'b0010101110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101110100100101101) && ({row_reg, col_reg}<22'b0010101110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101110101101010111) && ({row_reg, col_reg}<22'b0010101110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010101110101110000010) && ({row_reg, col_reg}<22'b0010101110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101110110000000010) && ({row_reg, col_reg}<22'b0010101110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101110110000101101) && ({row_reg, col_reg}<22'b0010101111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101111000001010111) && ({row_reg, col_reg}<22'b0010101111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101111000010000010) && ({row_reg, col_reg}<22'b0010101111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101111000100000010) && ({row_reg, col_reg}<22'b0010101111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101111000100101101) && ({row_reg, col_reg}<22'b0010101111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101111001101010111) && ({row_reg, col_reg}<22'b0010101111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010101111001110000010) && ({row_reg, col_reg}<22'b0010101111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101111010000000010) && ({row_reg, col_reg}<22'b0010101111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101111010000101101) && ({row_reg, col_reg}<22'b0010101111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101111100001010111) && ({row_reg, col_reg}<22'b0010101111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010101111100010000010) && ({row_reg, col_reg}<22'b0010101111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101111100100000010) && ({row_reg, col_reg}<22'b0010101111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101111100100101101) && ({row_reg, col_reg}<22'b0010101111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010101111101101010111) && ({row_reg, col_reg}<22'b0010101111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010101111101110000010) && ({row_reg, col_reg}<22'b0010101111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010101111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010101111110000000010) && ({row_reg, col_reg}<22'b0010101111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010101111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010101111110000101101) && ({row_reg, col_reg}<22'b0010110000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110000000001010111) && ({row_reg, col_reg}<22'b0010110000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110000000010000010) && ({row_reg, col_reg}<22'b0010110000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110000000100000010) && ({row_reg, col_reg}<22'b0010110000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110000000100101101) && ({row_reg, col_reg}<22'b0010110000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110000001101010111) && ({row_reg, col_reg}<22'b0010110000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010110000001110000010) && ({row_reg, col_reg}<22'b0010110000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110000010000000010) && ({row_reg, col_reg}<22'b0010110000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110000010000101101) && ({row_reg, col_reg}<22'b0010110000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110000100001010111) && ({row_reg, col_reg}<22'b0010110000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110000100010000010) && ({row_reg, col_reg}<22'b0010110000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110000100100000010) && ({row_reg, col_reg}<22'b0010110000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110000100100101101) && ({row_reg, col_reg}<22'b0010110000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110000101101010111) && ({row_reg, col_reg}<22'b0010110000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010110000101110000010) && ({row_reg, col_reg}<22'b0010110000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110000110000000010) && ({row_reg, col_reg}<22'b0010110000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110000110000101101) && ({row_reg, col_reg}<22'b0010110001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110001000001010111) && ({row_reg, col_reg}<22'b0010110001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110001000010000010) && ({row_reg, col_reg}<22'b0010110001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110001000100000010) && ({row_reg, col_reg}<22'b0010110001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110001000100101101) && ({row_reg, col_reg}<22'b0010110001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110001001101010111) && ({row_reg, col_reg}<22'b0010110001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010110001001110000010) && ({row_reg, col_reg}<22'b0010110001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110001010000000010) && ({row_reg, col_reg}<22'b0010110001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110001010000101101) && ({row_reg, col_reg}<22'b0010110001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110001100001010111) && ({row_reg, col_reg}<22'b0010110001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110001100010000010) && ({row_reg, col_reg}<22'b0010110001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110001100100000010) && ({row_reg, col_reg}<22'b0010110001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110001100100101101) && ({row_reg, col_reg}<22'b0010110001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110001101101010111) && ({row_reg, col_reg}<22'b0010110001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110001101110000010) && ({row_reg, col_reg}<22'b0010110001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110001110000000010) && ({row_reg, col_reg}<22'b0010110001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110001110000101101) && ({row_reg, col_reg}<22'b0010110010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110010000001010111) && ({row_reg, col_reg}<22'b0010110010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010110010000010000010) && ({row_reg, col_reg}<22'b0010110010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110010000100000010) && ({row_reg, col_reg}<22'b0010110010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110010000100101101) && ({row_reg, col_reg}<22'b0010110010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110010001101010111) && ({row_reg, col_reg}<22'b0010110010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110010001110000010) && ({row_reg, col_reg}<22'b0010110010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110010010000000010) && ({row_reg, col_reg}<22'b0010110010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110010010000101101) && ({row_reg, col_reg}<22'b0010110010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110010100001010111) && ({row_reg, col_reg}<22'b0010110010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010110010100010000010) && ({row_reg, col_reg}<22'b0010110010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110010100100000010) && ({row_reg, col_reg}<22'b0010110010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110010100100101101) && ({row_reg, col_reg}<22'b0010110010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110010101101010111) && ({row_reg, col_reg}<22'b0010110010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110010101110000010) && ({row_reg, col_reg}<22'b0010110010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110010110000000010) && ({row_reg, col_reg}<22'b0010110010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110010110000101101) && ({row_reg, col_reg}<22'b0010110011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110011000001010111) && ({row_reg, col_reg}<22'b0010110011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010110011000010000010) && ({row_reg, col_reg}<22'b0010110011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110011000100000010) && ({row_reg, col_reg}<22'b0010110011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110011000100101101) && ({row_reg, col_reg}<22'b0010110011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110011001101010111) && ({row_reg, col_reg}<22'b0010110011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110011001110000010) && ({row_reg, col_reg}<22'b0010110011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110011010000000010) && ({row_reg, col_reg}<22'b0010110011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110011010000101101) && ({row_reg, col_reg}<22'b0010110011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110011100001010111) && ({row_reg, col_reg}<22'b0010110011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010110011100010000010) && ({row_reg, col_reg}<22'b0010110011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110011100100000010) && ({row_reg, col_reg}<22'b0010110011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110011100100101101) && ({row_reg, col_reg}<22'b0010110011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110011101101010111) && ({row_reg, col_reg}<22'b0010110011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110011101110000010) && ({row_reg, col_reg}<22'b0010110011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110011110000000010) && ({row_reg, col_reg}<22'b0010110011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110011110000101101) && ({row_reg, col_reg}<22'b0010110100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110100000001010111) && ({row_reg, col_reg}<22'b0010110100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010110100000010000010) && ({row_reg, col_reg}<22'b0010110100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110100000100000010) && ({row_reg, col_reg}<22'b0010110100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110100000100101101) && ({row_reg, col_reg}<22'b0010110100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110100001101010111) && ({row_reg, col_reg}<22'b0010110100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110100001110000010) && ({row_reg, col_reg}<22'b0010110100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110100010000000010) && ({row_reg, col_reg}<22'b0010110100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110100010000101101) && ({row_reg, col_reg}<22'b0010110100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110100100001010111) && ({row_reg, col_reg}<22'b0010110100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010110100100010000010) && ({row_reg, col_reg}<22'b0010110100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110100100100000010) && ({row_reg, col_reg}<22'b0010110100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110100100100101101) && ({row_reg, col_reg}<22'b0010110100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110100101101010111) && ({row_reg, col_reg}<22'b0010110100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110100101110000010) && ({row_reg, col_reg}<22'b0010110100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110100110000000010) && ({row_reg, col_reg}<22'b0010110100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110100110000101101) && ({row_reg, col_reg}<22'b0010110101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110101000001010111) && ({row_reg, col_reg}<22'b0010110101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010110101000010000010) && ({row_reg, col_reg}<22'b0010110101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110101000100000010) && ({row_reg, col_reg}<22'b0010110101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110101000100101101) && ({row_reg, col_reg}<22'b0010110101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110101001101010111) && ({row_reg, col_reg}<22'b0010110101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110101001110000010) && ({row_reg, col_reg}<22'b0010110101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110101010000000010) && ({row_reg, col_reg}<22'b0010110101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110101010000101101) && ({row_reg, col_reg}<22'b0010110101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110101100001010111) && ({row_reg, col_reg}<22'b0010110101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110101100010000010) && ({row_reg, col_reg}<22'b0010110101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110101100100000010) && ({row_reg, col_reg}<22'b0010110101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110101100100101101) && ({row_reg, col_reg}<22'b0010110101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110101101101010111) && ({row_reg, col_reg}<22'b0010110101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110101101110000010) && ({row_reg, col_reg}<22'b0010110101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110101110000000010) && ({row_reg, col_reg}<22'b0010110101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110101110000101101) && ({row_reg, col_reg}<22'b0010110110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110110000001010111) && ({row_reg, col_reg}<22'b0010110110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110110000010000010) && ({row_reg, col_reg}<22'b0010110110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110110000100000010) && ({row_reg, col_reg}<22'b0010110110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110110000100101101) && ({row_reg, col_reg}<22'b0010110110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110110001101010111) && ({row_reg, col_reg}<22'b0010110110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110110001110000010) && ({row_reg, col_reg}<22'b0010110110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110110010000000010) && ({row_reg, col_reg}<22'b0010110110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110110010000101101) && ({row_reg, col_reg}<22'b0010110110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110110100001010111) && ({row_reg, col_reg}<22'b0010110110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110110100010000010) && ({row_reg, col_reg}<22'b0010110110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110110100100000010) && ({row_reg, col_reg}<22'b0010110110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110110100100101101) && ({row_reg, col_reg}<22'b0010110110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110110101101010111) && ({row_reg, col_reg}<22'b0010110110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110110101110000010) && ({row_reg, col_reg}<22'b0010110110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110110110000000010) && ({row_reg, col_reg}<22'b0010110110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110110110000101101) && ({row_reg, col_reg}<22'b0010110111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110111000001010111) && ({row_reg, col_reg}<22'b0010110111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110111000010000010) && ({row_reg, col_reg}<22'b0010110111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110111000100000010) && ({row_reg, col_reg}<22'b0010110111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110111000100101101) && ({row_reg, col_reg}<22'b0010110111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110111001101010111) && ({row_reg, col_reg}<22'b0010110111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110111001110000010) && ({row_reg, col_reg}<22'b0010110111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110111010000000010) && ({row_reg, col_reg}<22'b0010110111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110111010000101101) && ({row_reg, col_reg}<22'b0010110111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110111100001010111) && ({row_reg, col_reg}<22'b0010110111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110111100010000010) && ({row_reg, col_reg}<22'b0010110111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110111100100000010) && ({row_reg, col_reg}<22'b0010110111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110111100100101101) && ({row_reg, col_reg}<22'b0010110111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010110111101101010111) && ({row_reg, col_reg}<22'b0010110111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010110111101110000010) && ({row_reg, col_reg}<22'b0010110111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010110111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010110111110000000010) && ({row_reg, col_reg}<22'b0010110111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010110111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010110111110000101101) && ({row_reg, col_reg}<22'b0010111000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111000000001010111) && ({row_reg, col_reg}<22'b0010111000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111000000010000010) && ({row_reg, col_reg}<22'b0010111000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111000000100000010) && ({row_reg, col_reg}<22'b0010111000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111000000100101101) && ({row_reg, col_reg}<22'b0010111000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111000001101010111) && ({row_reg, col_reg}<22'b0010111000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111000001110000010) && ({row_reg, col_reg}<22'b0010111000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111000010000000010) && ({row_reg, col_reg}<22'b0010111000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111000010000101101) && ({row_reg, col_reg}<22'b0010111000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111000100001010111) && ({row_reg, col_reg}<22'b0010111000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111000100010000010) && ({row_reg, col_reg}<22'b0010111000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111000100100000010) && ({row_reg, col_reg}<22'b0010111000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111000100100101101) && ({row_reg, col_reg}<22'b0010111000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111000101101010111) && ({row_reg, col_reg}<22'b0010111000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111000101110000010) && ({row_reg, col_reg}<22'b0010111000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111000110000000010) && ({row_reg, col_reg}<22'b0010111000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111000110000101101) && ({row_reg, col_reg}<22'b0010111001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111001000001010111) && ({row_reg, col_reg}<22'b0010111001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111001000010000010) && ({row_reg, col_reg}<22'b0010111001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111001000100000010) && ({row_reg, col_reg}<22'b0010111001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111001000100101101) && ({row_reg, col_reg}<22'b0010111001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111001001101010111) && ({row_reg, col_reg}<22'b0010111001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010111001001110000010) && ({row_reg, col_reg}<22'b0010111001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111001010000000010) && ({row_reg, col_reg}<22'b0010111001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111001010000101101) && ({row_reg, col_reg}<22'b0010111001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111001100001010111) && ({row_reg, col_reg}<22'b0010111001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111001100010000010) && ({row_reg, col_reg}<22'b0010111001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111001100100000010) && ({row_reg, col_reg}<22'b0010111001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111001100100101101) && ({row_reg, col_reg}<22'b0010111001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111001101101010111) && ({row_reg, col_reg}<22'b0010111001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010111001101110000010) && ({row_reg, col_reg}<22'b0010111001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111001110000000010) && ({row_reg, col_reg}<22'b0010111001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111001110000101101) && ({row_reg, col_reg}<22'b0010111010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111010000001010111) && ({row_reg, col_reg}<22'b0010111010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111010000010000010) && ({row_reg, col_reg}<22'b0010111010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111010000100000010) && ({row_reg, col_reg}<22'b0010111010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111010000100101101) && ({row_reg, col_reg}<22'b0010111010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111010001101010111) && ({row_reg, col_reg}<22'b0010111010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010111010001110000010) && ({row_reg, col_reg}<22'b0010111010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111010010000000010) && ({row_reg, col_reg}<22'b0010111010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111010010000101101) && ({row_reg, col_reg}<22'b0010111010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111010100001010111) && ({row_reg, col_reg}<22'b0010111010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111010100010000010) && ({row_reg, col_reg}<22'b0010111010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111010100100000010) && ({row_reg, col_reg}<22'b0010111010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111010100100101101) && ({row_reg, col_reg}<22'b0010111010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111010101101010111) && ({row_reg, col_reg}<22'b0010111010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111010101110000010) && ({row_reg, col_reg}<22'b0010111010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111010110000000010) && ({row_reg, col_reg}<22'b0010111010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111010110000101101) && ({row_reg, col_reg}<22'b0010111011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111011000001010111) && ({row_reg, col_reg}<22'b0010111011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111011000010000010) && ({row_reg, col_reg}<22'b0010111011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111011000100000010) && ({row_reg, col_reg}<22'b0010111011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111011000100101101) && ({row_reg, col_reg}<22'b0010111011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111011001101010111) && ({row_reg, col_reg}<22'b0010111011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111011001110000010) && ({row_reg, col_reg}<22'b0010111011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111011010000000010) && ({row_reg, col_reg}<22'b0010111011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111011010000101101) && ({row_reg, col_reg}<22'b0010111011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111011100001010111) && ({row_reg, col_reg}<22'b0010111011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111011100010000010) && ({row_reg, col_reg}<22'b0010111011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111011100100000010) && ({row_reg, col_reg}<22'b0010111011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111011100100101101) && ({row_reg, col_reg}<22'b0010111011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111011101101010111) && ({row_reg, col_reg}<22'b0010111011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111011101110000010) && ({row_reg, col_reg}<22'b0010111011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111011110000000010) && ({row_reg, col_reg}<22'b0010111011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111011110000101101) && ({row_reg, col_reg}<22'b0010111100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111100000001010111) && ({row_reg, col_reg}<22'b0010111100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111100000010000010) && ({row_reg, col_reg}<22'b0010111100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111100000100000010) && ({row_reg, col_reg}<22'b0010111100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111100000100101101) && ({row_reg, col_reg}<22'b0010111100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111100001101010111) && ({row_reg, col_reg}<22'b0010111100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111100001110000010) && ({row_reg, col_reg}<22'b0010111100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111100010000000010) && ({row_reg, col_reg}<22'b0010111100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111100010000101101) && ({row_reg, col_reg}<22'b0010111100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111100100001010111) && ({row_reg, col_reg}<22'b0010111100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111100100010000010) && ({row_reg, col_reg}<22'b0010111100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111100100100000010) && ({row_reg, col_reg}<22'b0010111100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111100100100101101) && ({row_reg, col_reg}<22'b0010111100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111100101101010111) && ({row_reg, col_reg}<22'b0010111100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111100101110000010) && ({row_reg, col_reg}<22'b0010111100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111100110000000010) && ({row_reg, col_reg}<22'b0010111100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111100110000101101) && ({row_reg, col_reg}<22'b0010111101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111101000001010111) && ({row_reg, col_reg}<22'b0010111101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010111101000010000010) && ({row_reg, col_reg}<22'b0010111101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111101000100000010) && ({row_reg, col_reg}<22'b0010111101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111101000100101101) && ({row_reg, col_reg}<22'b0010111101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111101001101010111) && ({row_reg, col_reg}<22'b0010111101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111101001110000010) && ({row_reg, col_reg}<22'b0010111101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111101010000000010) && ({row_reg, col_reg}<22'b0010111101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111101010000101101) && ({row_reg, col_reg}<22'b0010111101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111101100001010111) && ({row_reg, col_reg}<22'b0010111101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010111101100010000010) && ({row_reg, col_reg}<22'b0010111101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111101100100000010) && ({row_reg, col_reg}<22'b0010111101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111101100100101101) && ({row_reg, col_reg}<22'b0010111101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111101101101010111) && ({row_reg, col_reg}<22'b0010111101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111101101110000010) && ({row_reg, col_reg}<22'b0010111101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111101110000000010) && ({row_reg, col_reg}<22'b0010111101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111101110000101101) && ({row_reg, col_reg}<22'b0010111110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111110000001010111) && ({row_reg, col_reg}<22'b0010111110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0010111110000010000010) && ({row_reg, col_reg}<22'b0010111110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111110000100000010) && ({row_reg, col_reg}<22'b0010111110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111110000100101101) && ({row_reg, col_reg}<22'b0010111110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111110001101010111) && ({row_reg, col_reg}<22'b0010111110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111110001110000010) && ({row_reg, col_reg}<22'b0010111110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111110010000000010) && ({row_reg, col_reg}<22'b0010111110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111110010000101101) && ({row_reg, col_reg}<22'b0010111110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111110100001010111) && ({row_reg, col_reg}<22'b0010111110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111110100010000010) && ({row_reg, col_reg}<22'b0010111110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111110100100000010) && ({row_reg, col_reg}<22'b0010111110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111110100100101101) && ({row_reg, col_reg}<22'b0010111110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111110101101010111) && ({row_reg, col_reg}<22'b0010111110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111110101110000010) && ({row_reg, col_reg}<22'b0010111110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111110110000000010) && ({row_reg, col_reg}<22'b0010111110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111110110000101101) && ({row_reg, col_reg}<22'b0010111111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111111000001010111) && ({row_reg, col_reg}<22'b0010111111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0010111111000010000010) && ({row_reg, col_reg}<22'b0010111111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111111000100000010) && ({row_reg, col_reg}<22'b0010111111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111111000100101101) && ({row_reg, col_reg}<22'b0010111111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111111001101010111) && ({row_reg, col_reg}<22'b0010111111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111111001110000010) && ({row_reg, col_reg}<22'b0010111111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111111010000000010) && ({row_reg, col_reg}<22'b0010111111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111111010000101101) && ({row_reg, col_reg}<22'b0010111111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111111100001010111) && ({row_reg, col_reg}<22'b0010111111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111111100010000010) && ({row_reg, col_reg}<22'b0010111111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111111100100000010) && ({row_reg, col_reg}<22'b0010111111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111111100100101101) && ({row_reg, col_reg}<22'b0010111111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0010111111101101010111) && ({row_reg, col_reg}<22'b0010111111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0010111111101110000010) && ({row_reg, col_reg}<22'b0010111111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0010111111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0010111111110000000010) && ({row_reg, col_reg}<22'b0010111111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0010111111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0010111111110000101101) && ({row_reg, col_reg}<22'b0011000000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000000000001010111) && ({row_reg, col_reg}<22'b0011000000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000000000010000010) && ({row_reg, col_reg}<22'b0011000000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000000000100000010) && ({row_reg, col_reg}<22'b0011000000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000000000100101101) && ({row_reg, col_reg}<22'b0011000000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000000001101010111) && ({row_reg, col_reg}<22'b0011000000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000000001110000010) && ({row_reg, col_reg}<22'b0011000000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000000010000000010) && ({row_reg, col_reg}<22'b0011000000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000000010000101101) && ({row_reg, col_reg}<22'b0011000000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000000100001010111) && ({row_reg, col_reg}<22'b0011000000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000000100010000010) && ({row_reg, col_reg}<22'b0011000000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000000100100000010) && ({row_reg, col_reg}<22'b0011000000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000000100100101101) && ({row_reg, col_reg}<22'b0011000000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000000101101010111) && ({row_reg, col_reg}<22'b0011000000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000000101110000010) && ({row_reg, col_reg}<22'b0011000000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000000110000000010) && ({row_reg, col_reg}<22'b0011000000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000000110000101101) && ({row_reg, col_reg}<22'b0011000001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000001000001010111) && ({row_reg, col_reg}<22'b0011000001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000001000010000010) && ({row_reg, col_reg}<22'b0011000001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000001000100000010) && ({row_reg, col_reg}<22'b0011000001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000001000100101101) && ({row_reg, col_reg}<22'b0011000001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000001001101010111) && ({row_reg, col_reg}<22'b0011000001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000001001110000010) && ({row_reg, col_reg}<22'b0011000001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000001010000000010) && ({row_reg, col_reg}<22'b0011000001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000001010000101101) && ({row_reg, col_reg}<22'b0011000001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000001100001010111) && ({row_reg, col_reg}<22'b0011000001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000001100010000010) && ({row_reg, col_reg}<22'b0011000001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000001100100000010) && ({row_reg, col_reg}<22'b0011000001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000001100100101101) && ({row_reg, col_reg}<22'b0011000001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000001101101010111) && ({row_reg, col_reg}<22'b0011000001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000001101110000010) && ({row_reg, col_reg}<22'b0011000001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000001110000000010) && ({row_reg, col_reg}<22'b0011000001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000001110000101101) && ({row_reg, col_reg}<22'b0011000010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000010000001010111) && ({row_reg, col_reg}<22'b0011000010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000010000010000010) && ({row_reg, col_reg}<22'b0011000010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000010000100000010) && ({row_reg, col_reg}<22'b0011000010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000010000100101101) && ({row_reg, col_reg}<22'b0011000010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000010001101010111) && ({row_reg, col_reg}<22'b0011000010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011000010001110000010) && ({row_reg, col_reg}<22'b0011000010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000010010000000010) && ({row_reg, col_reg}<22'b0011000010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000010010000101101) && ({row_reg, col_reg}<22'b0011000010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000010100001010111) && ({row_reg, col_reg}<22'b0011000010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000010100010000010) && ({row_reg, col_reg}<22'b0011000010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000010100100000010) && ({row_reg, col_reg}<22'b0011000010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000010100100101101) && ({row_reg, col_reg}<22'b0011000010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000010101101010111) && ({row_reg, col_reg}<22'b0011000010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011000010101110000010) && ({row_reg, col_reg}<22'b0011000010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000010110000000010) && ({row_reg, col_reg}<22'b0011000010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000010110000101101) && ({row_reg, col_reg}<22'b0011000011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000011000001010111) && ({row_reg, col_reg}<22'b0011000011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000011000010000010) && ({row_reg, col_reg}<22'b0011000011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000011000100000010) && ({row_reg, col_reg}<22'b0011000011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000011000100101101) && ({row_reg, col_reg}<22'b0011000011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000011001101010111) && ({row_reg, col_reg}<22'b0011000011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011000011001110000010) && ({row_reg, col_reg}<22'b0011000011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000011010000000010) && ({row_reg, col_reg}<22'b0011000011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000011010000101101) && ({row_reg, col_reg}<22'b0011000011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000011100001010111) && ({row_reg, col_reg}<22'b0011000011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000011100010000010) && ({row_reg, col_reg}<22'b0011000011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000011100100000010) && ({row_reg, col_reg}<22'b0011000011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000011100100101101) && ({row_reg, col_reg}<22'b0011000011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000011101101010111) && ({row_reg, col_reg}<22'b0011000011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011000011101110000010) && ({row_reg, col_reg}<22'b0011000011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000011110000000010) && ({row_reg, col_reg}<22'b0011000011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000011110000101101) && ({row_reg, col_reg}<22'b0011000100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000100000001010111) && ({row_reg, col_reg}<22'b0011000100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000100000010000010) && ({row_reg, col_reg}<22'b0011000100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000100000100000010) && ({row_reg, col_reg}<22'b0011000100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000100000100101101) && ({row_reg, col_reg}<22'b0011000100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000100001101010111) && ({row_reg, col_reg}<22'b0011000100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011000100001110000010) && ({row_reg, col_reg}<22'b0011000100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000100010000000010) && ({row_reg, col_reg}<22'b0011000100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000100010000101101) && ({row_reg, col_reg}<22'b0011000100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000100100001010111) && ({row_reg, col_reg}<22'b0011000100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000100100010000010) && ({row_reg, col_reg}<22'b0011000100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000100100100000010) && ({row_reg, col_reg}<22'b0011000100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000100100100101101) && ({row_reg, col_reg}<22'b0011000100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000100101101010111) && ({row_reg, col_reg}<22'b0011000100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011000100101110000010) && ({row_reg, col_reg}<22'b0011000100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000100110000000010) && ({row_reg, col_reg}<22'b0011000100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000100110000101101) && ({row_reg, col_reg}<22'b0011000101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000101000001010111) && ({row_reg, col_reg}<22'b0011000101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000101000010000010) && ({row_reg, col_reg}<22'b0011000101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000101000100000010) && ({row_reg, col_reg}<22'b0011000101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000101000100101101) && ({row_reg, col_reg}<22'b0011000101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000101001101010111) && ({row_reg, col_reg}<22'b0011000101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011000101001110000010) && ({row_reg, col_reg}<22'b0011000101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000101010000000010) && ({row_reg, col_reg}<22'b0011000101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000101010000101101) && ({row_reg, col_reg}<22'b0011000101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000101100001010111) && ({row_reg, col_reg}<22'b0011000101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000101100010000010) && ({row_reg, col_reg}<22'b0011000101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000101100100000010) && ({row_reg, col_reg}<22'b0011000101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000101100100101101) && ({row_reg, col_reg}<22'b0011000101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000101101101010111) && ({row_reg, col_reg}<22'b0011000101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000101101110000010) && ({row_reg, col_reg}<22'b0011000101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000101110000000010) && ({row_reg, col_reg}<22'b0011000101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000101110000101101) && ({row_reg, col_reg}<22'b0011000110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000110000001010111) && ({row_reg, col_reg}<22'b0011000110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011000110000010000010) && ({row_reg, col_reg}<22'b0011000110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000110000100000010) && ({row_reg, col_reg}<22'b0011000110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000110000100101101) && ({row_reg, col_reg}<22'b0011000110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000110001101010111) && ({row_reg, col_reg}<22'b0011000110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000110001110000010) && ({row_reg, col_reg}<22'b0011000110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000110010000000010) && ({row_reg, col_reg}<22'b0011000110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000110010000101101) && ({row_reg, col_reg}<22'b0011000110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000110100001010111) && ({row_reg, col_reg}<22'b0011000110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011000110100010000010) && ({row_reg, col_reg}<22'b0011000110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000110100100000010) && ({row_reg, col_reg}<22'b0011000110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000110100100101101) && ({row_reg, col_reg}<22'b0011000110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000110101101010111) && ({row_reg, col_reg}<22'b0011000110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000110101110000010) && ({row_reg, col_reg}<22'b0011000110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000110110000000010) && ({row_reg, col_reg}<22'b0011000110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000110110000101101) && ({row_reg, col_reg}<22'b0011000111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000111000001010111) && ({row_reg, col_reg}<22'b0011000111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011000111000010000010) && ({row_reg, col_reg}<22'b0011000111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000111000100000010) && ({row_reg, col_reg}<22'b0011000111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000111000100101101) && ({row_reg, col_reg}<22'b0011000111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000111001101010111) && ({row_reg, col_reg}<22'b0011000111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000111001110000010) && ({row_reg, col_reg}<22'b0011000111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000111010000000010) && ({row_reg, col_reg}<22'b0011000111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000111010000101101) && ({row_reg, col_reg}<22'b0011000111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000111100001010111) && ({row_reg, col_reg}<22'b0011000111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011000111100010000010) && ({row_reg, col_reg}<22'b0011000111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000111100100000010) && ({row_reg, col_reg}<22'b0011000111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000111100100101101) && ({row_reg, col_reg}<22'b0011000111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011000111101101010111) && ({row_reg, col_reg}<22'b0011000111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011000111101110000010) && ({row_reg, col_reg}<22'b0011000111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011000111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011000111110000000010) && ({row_reg, col_reg}<22'b0011000111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011000111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011000111110000101101) && ({row_reg, col_reg}<22'b0011001000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001000000001010111) && ({row_reg, col_reg}<22'b0011001000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011001000000010000010) && ({row_reg, col_reg}<22'b0011001000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001000000100000010) && ({row_reg, col_reg}<22'b0011001000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001000000100101101) && ({row_reg, col_reg}<22'b0011001000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001000001101010111) && ({row_reg, col_reg}<22'b0011001000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001000001110000010) && ({row_reg, col_reg}<22'b0011001000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001000010000000010) && ({row_reg, col_reg}<22'b0011001000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001000010000101101) && ({row_reg, col_reg}<22'b0011001000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001000100001010111) && ({row_reg, col_reg}<22'b0011001000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011001000100010000010) && ({row_reg, col_reg}<22'b0011001000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001000100100000010) && ({row_reg, col_reg}<22'b0011001000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001000100100101101) && ({row_reg, col_reg}<22'b0011001000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001000101101010111) && ({row_reg, col_reg}<22'b0011001000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001000101110000010) && ({row_reg, col_reg}<22'b0011001000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001000110000000010) && ({row_reg, col_reg}<22'b0011001000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001000110000101101) && ({row_reg, col_reg}<22'b0011001001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001001000001010111) && ({row_reg, col_reg}<22'b0011001001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011001001000010000010) && ({row_reg, col_reg}<22'b0011001001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001001000100000010) && ({row_reg, col_reg}<22'b0011001001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001001000100101101) && ({row_reg, col_reg}<22'b0011001001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001001001101010111) && ({row_reg, col_reg}<22'b0011001001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001001001110000010) && ({row_reg, col_reg}<22'b0011001001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001001010000000010) && ({row_reg, col_reg}<22'b0011001001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001001010000101101) && ({row_reg, col_reg}<22'b0011001001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001001100001010111) && ({row_reg, col_reg}<22'b0011001001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001001100010000010) && ({row_reg, col_reg}<22'b0011001001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001001100100000010) && ({row_reg, col_reg}<22'b0011001001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001001100100101101) && ({row_reg, col_reg}<22'b0011001001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001001101101010111) && ({row_reg, col_reg}<22'b0011001001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001001101110000010) && ({row_reg, col_reg}<22'b0011001001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001001110000000010) && ({row_reg, col_reg}<22'b0011001001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001001110000101101) && ({row_reg, col_reg}<22'b0011001010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001010000001010111) && ({row_reg, col_reg}<22'b0011001010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001010000010000010) && ({row_reg, col_reg}<22'b0011001010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001010000100000010) && ({row_reg, col_reg}<22'b0011001010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001010000100101101) && ({row_reg, col_reg}<22'b0011001010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001010001101010111) && ({row_reg, col_reg}<22'b0011001010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001010001110000010) && ({row_reg, col_reg}<22'b0011001010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001010010000000010) && ({row_reg, col_reg}<22'b0011001010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001010010000101101) && ({row_reg, col_reg}<22'b0011001010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001010100001010111) && ({row_reg, col_reg}<22'b0011001010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001010100010000010) && ({row_reg, col_reg}<22'b0011001010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001010100100000010) && ({row_reg, col_reg}<22'b0011001010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001010100100101101) && ({row_reg, col_reg}<22'b0011001010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001010101101010111) && ({row_reg, col_reg}<22'b0011001010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001010101110000010) && ({row_reg, col_reg}<22'b0011001010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001010110000000010) && ({row_reg, col_reg}<22'b0011001010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001010110000101101) && ({row_reg, col_reg}<22'b0011001011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001011000001010111) && ({row_reg, col_reg}<22'b0011001011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001011000010000010) && ({row_reg, col_reg}<22'b0011001011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001011000100000010) && ({row_reg, col_reg}<22'b0011001011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001011000100101101) && ({row_reg, col_reg}<22'b0011001011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001011001101010111) && ({row_reg, col_reg}<22'b0011001011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001011001110000010) && ({row_reg, col_reg}<22'b0011001011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001011010000000010) && ({row_reg, col_reg}<22'b0011001011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001011010000101101) && ({row_reg, col_reg}<22'b0011001011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001011100001010111) && ({row_reg, col_reg}<22'b0011001011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001011100010000010) && ({row_reg, col_reg}<22'b0011001011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001011100100000010) && ({row_reg, col_reg}<22'b0011001011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001011100100101101) && ({row_reg, col_reg}<22'b0011001011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001011101101010111) && ({row_reg, col_reg}<22'b0011001011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001011101110000010) && ({row_reg, col_reg}<22'b0011001011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001011110000000010) && ({row_reg, col_reg}<22'b0011001011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001011110000101101) && ({row_reg, col_reg}<22'b0011001100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001100000001010111) && ({row_reg, col_reg}<22'b0011001100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001100000010000010) && ({row_reg, col_reg}<22'b0011001100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001100000100000010) && ({row_reg, col_reg}<22'b0011001100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001100000100101101) && ({row_reg, col_reg}<22'b0011001100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001100001101010111) && ({row_reg, col_reg}<22'b0011001100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011001100001110000010) && ({row_reg, col_reg}<22'b0011001100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001100010000000010) && ({row_reg, col_reg}<22'b0011001100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001100010000101101) && ({row_reg, col_reg}<22'b0011001100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001100100001010111) && ({row_reg, col_reg}<22'b0011001100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001100100010000010) && ({row_reg, col_reg}<22'b0011001100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001100100100000010) && ({row_reg, col_reg}<22'b0011001100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001100100100101101) && ({row_reg, col_reg}<22'b0011001100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001100101101010111) && ({row_reg, col_reg}<22'b0011001100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011001100101110000010) && ({row_reg, col_reg}<22'b0011001100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001100110000000010) && ({row_reg, col_reg}<22'b0011001100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001100110000101101) && ({row_reg, col_reg}<22'b0011001101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001101000001010111) && ({row_reg, col_reg}<22'b0011001101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001101000010000010) && ({row_reg, col_reg}<22'b0011001101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001101000100000010) && ({row_reg, col_reg}<22'b0011001101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001101000100101101) && ({row_reg, col_reg}<22'b0011001101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001101001101010111) && ({row_reg, col_reg}<22'b0011001101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011001101001110000010) && ({row_reg, col_reg}<22'b0011001101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001101010000000010) && ({row_reg, col_reg}<22'b0011001101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001101010000101101) && ({row_reg, col_reg}<22'b0011001101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001101100001010111) && ({row_reg, col_reg}<22'b0011001101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001101100010000010) && ({row_reg, col_reg}<22'b0011001101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001101100100000010) && ({row_reg, col_reg}<22'b0011001101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001101100100101101) && ({row_reg, col_reg}<22'b0011001101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001101101101010111) && ({row_reg, col_reg}<22'b0011001101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011001101101110000010) && ({row_reg, col_reg}<22'b0011001101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001101110000000010) && ({row_reg, col_reg}<22'b0011001101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001101110000101101) && ({row_reg, col_reg}<22'b0011001110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001110000001010111) && ({row_reg, col_reg}<22'b0011001110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001110000010000010) && ({row_reg, col_reg}<22'b0011001110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001110000100000010) && ({row_reg, col_reg}<22'b0011001110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001110000100101101) && ({row_reg, col_reg}<22'b0011001110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001110001101010111) && ({row_reg, col_reg}<22'b0011001110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011001110001110000010) && ({row_reg, col_reg}<22'b0011001110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001110010000000010) && ({row_reg, col_reg}<22'b0011001110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001110010000101101) && ({row_reg, col_reg}<22'b0011001110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001110100001010111) && ({row_reg, col_reg}<22'b0011001110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001110100010000010) && ({row_reg, col_reg}<22'b0011001110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001110100100000010) && ({row_reg, col_reg}<22'b0011001110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001110100100101101) && ({row_reg, col_reg}<22'b0011001110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001110101101010111) && ({row_reg, col_reg}<22'b0011001110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011001110101110000010) && ({row_reg, col_reg}<22'b0011001110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001110110000000010) && ({row_reg, col_reg}<22'b0011001110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001110110000101101) && ({row_reg, col_reg}<22'b0011001111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001111000001010111) && ({row_reg, col_reg}<22'b0011001111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001111000010000010) && ({row_reg, col_reg}<22'b0011001111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001111000100000010) && ({row_reg, col_reg}<22'b0011001111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001111000100101101) && ({row_reg, col_reg}<22'b0011001111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001111001101010111) && ({row_reg, col_reg}<22'b0011001111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011001111001110000010) && ({row_reg, col_reg}<22'b0011001111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001111010000000010) && ({row_reg, col_reg}<22'b0011001111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001111010000101101) && ({row_reg, col_reg}<22'b0011001111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001111100001010111) && ({row_reg, col_reg}<22'b0011001111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001111100010000010) && ({row_reg, col_reg}<22'b0011001111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001111100100000010) && ({row_reg, col_reg}<22'b0011001111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001111100100101101) && ({row_reg, col_reg}<22'b0011001111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011001111101101010111) && ({row_reg, col_reg}<22'b0011001111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011001111101110000010) && ({row_reg, col_reg}<22'b0011001111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011001111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011001111110000000010) && ({row_reg, col_reg}<22'b0011001111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011001111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011001111110000101101) && ({row_reg, col_reg}<22'b0011010000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010000000001010111) && ({row_reg, col_reg}<22'b0011010000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011010000000010000010) && ({row_reg, col_reg}<22'b0011010000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010000000100000010) && ({row_reg, col_reg}<22'b0011010000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010000000100101101) && ({row_reg, col_reg}<22'b0011010000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010000001101010111) && ({row_reg, col_reg}<22'b0011010000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010000001110000010) && ({row_reg, col_reg}<22'b0011010000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010000010000000010) && ({row_reg, col_reg}<22'b0011010000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010000010000101101) && ({row_reg, col_reg}<22'b0011010000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010000100001010111) && ({row_reg, col_reg}<22'b0011010000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011010000100010000010) && ({row_reg, col_reg}<22'b0011010000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010000100100000010) && ({row_reg, col_reg}<22'b0011010000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010000100100101101) && ({row_reg, col_reg}<22'b0011010000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010000101101010111) && ({row_reg, col_reg}<22'b0011010000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010000101110000010) && ({row_reg, col_reg}<22'b0011010000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010000110000000010) && ({row_reg, col_reg}<22'b0011010000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010000110000101101) && ({row_reg, col_reg}<22'b0011010001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010001000001010111) && ({row_reg, col_reg}<22'b0011010001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011010001000010000010) && ({row_reg, col_reg}<22'b0011010001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010001000100000010) && ({row_reg, col_reg}<22'b0011010001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010001000100101101) && ({row_reg, col_reg}<22'b0011010001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010001001101010111) && ({row_reg, col_reg}<22'b0011010001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010001001110000010) && ({row_reg, col_reg}<22'b0011010001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010001010000000010) && ({row_reg, col_reg}<22'b0011010001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010001010000101101) && ({row_reg, col_reg}<22'b0011010001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010001100001010111) && ({row_reg, col_reg}<22'b0011010001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011010001100010000010) && ({row_reg, col_reg}<22'b0011010001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010001100100000010) && ({row_reg, col_reg}<22'b0011010001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010001100100101101) && ({row_reg, col_reg}<22'b0011010001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010001101101010111) && ({row_reg, col_reg}<22'b0011010001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010001101110000010) && ({row_reg, col_reg}<22'b0011010001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010001110000000010) && ({row_reg, col_reg}<22'b0011010001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010001110000101101) && ({row_reg, col_reg}<22'b0011010010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010010000001010111) && ({row_reg, col_reg}<22'b0011010010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011010010000010000010) && ({row_reg, col_reg}<22'b0011010010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010010000100000010) && ({row_reg, col_reg}<22'b0011010010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010010000100101101) && ({row_reg, col_reg}<22'b0011010010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010010001101010111) && ({row_reg, col_reg}<22'b0011010010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010010001110000010) && ({row_reg, col_reg}<22'b0011010010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010010010000000010) && ({row_reg, col_reg}<22'b0011010010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010010010000101101) && ({row_reg, col_reg}<22'b0011010010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010010100001010111) && ({row_reg, col_reg}<22'b0011010010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011010010100010000010) && ({row_reg, col_reg}<22'b0011010010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010010100100000010) && ({row_reg, col_reg}<22'b0011010010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010010100100101101) && ({row_reg, col_reg}<22'b0011010010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010010101101010111) && ({row_reg, col_reg}<22'b0011010010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010010101110000010) && ({row_reg, col_reg}<22'b0011010010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010010110000000010) && ({row_reg, col_reg}<22'b0011010010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010010110000101101) && ({row_reg, col_reg}<22'b0011010011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010011000001010111) && ({row_reg, col_reg}<22'b0011010011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011010011000010000010) && ({row_reg, col_reg}<22'b0011010011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010011000100000010) && ({row_reg, col_reg}<22'b0011010011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010011000100101101) && ({row_reg, col_reg}<22'b0011010011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010011001101010111) && ({row_reg, col_reg}<22'b0011010011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010011001110000010) && ({row_reg, col_reg}<22'b0011010011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010011010000000010) && ({row_reg, col_reg}<22'b0011010011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010011010000101101) && ({row_reg, col_reg}<22'b0011010011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010011100001010111) && ({row_reg, col_reg}<22'b0011010011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010011100010000010) && ({row_reg, col_reg}<22'b0011010011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010011100100000010) && ({row_reg, col_reg}<22'b0011010011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010011100100101101) && ({row_reg, col_reg}<22'b0011010011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010011101101010111) && ({row_reg, col_reg}<22'b0011010011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010011101110000010) && ({row_reg, col_reg}<22'b0011010011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010011110000000010) && ({row_reg, col_reg}<22'b0011010011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010011110000101101) && ({row_reg, col_reg}<22'b0011010100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010100000001010111) && ({row_reg, col_reg}<22'b0011010100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010100000010000010) && ({row_reg, col_reg}<22'b0011010100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010100000100000010) && ({row_reg, col_reg}<22'b0011010100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010100000100101101) && ({row_reg, col_reg}<22'b0011010100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010100001101010111) && ({row_reg, col_reg}<22'b0011010100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010100001110000010) && ({row_reg, col_reg}<22'b0011010100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010100010000000010) && ({row_reg, col_reg}<22'b0011010100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010100010000101101) && ({row_reg, col_reg}<22'b0011010100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010100100001010111) && ({row_reg, col_reg}<22'b0011010100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010100100010000010) && ({row_reg, col_reg}<22'b0011010100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010100100100000010) && ({row_reg, col_reg}<22'b0011010100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010100100100101101) && ({row_reg, col_reg}<22'b0011010100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010100101101010111) && ({row_reg, col_reg}<22'b0011010100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010100101110000010) && ({row_reg, col_reg}<22'b0011010100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010100110000000010) && ({row_reg, col_reg}<22'b0011010100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010100110000101101) && ({row_reg, col_reg}<22'b0011010101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010101000001010111) && ({row_reg, col_reg}<22'b0011010101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010101000010000010) && ({row_reg, col_reg}<22'b0011010101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010101000100000010) && ({row_reg, col_reg}<22'b0011010101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010101000100101101) && ({row_reg, col_reg}<22'b0011010101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010101001101010111) && ({row_reg, col_reg}<22'b0011010101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010101001110000010) && ({row_reg, col_reg}<22'b0011010101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010101010000000010) && ({row_reg, col_reg}<22'b0011010101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010101010000101101) && ({row_reg, col_reg}<22'b0011010101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010101100001010111) && ({row_reg, col_reg}<22'b0011010101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010101100010000010) && ({row_reg, col_reg}<22'b0011010101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010101100100000010) && ({row_reg, col_reg}<22'b0011010101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010101100100101101) && ({row_reg, col_reg}<22'b0011010101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010101101101010111) && ({row_reg, col_reg}<22'b0011010101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010101101110000010) && ({row_reg, col_reg}<22'b0011010101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010101110000000010) && ({row_reg, col_reg}<22'b0011010101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010101110000101101) && ({row_reg, col_reg}<22'b0011010110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010110000001010111) && ({row_reg, col_reg}<22'b0011010110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010110000010000010) && ({row_reg, col_reg}<22'b0011010110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010110000100000010) && ({row_reg, col_reg}<22'b0011010110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010110000100101101) && ({row_reg, col_reg}<22'b0011010110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010110001101010111) && ({row_reg, col_reg}<22'b0011010110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011010110001110000010) && ({row_reg, col_reg}<22'b0011010110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010110010000000010) && ({row_reg, col_reg}<22'b0011010110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010110010000101101) && ({row_reg, col_reg}<22'b0011010110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010110100001010111) && ({row_reg, col_reg}<22'b0011010110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010110100010000010) && ({row_reg, col_reg}<22'b0011010110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010110100100000010) && ({row_reg, col_reg}<22'b0011010110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010110100100101101) && ({row_reg, col_reg}<22'b0011010110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010110101101010111) && ({row_reg, col_reg}<22'b0011010110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011010110101110000010) && ({row_reg, col_reg}<22'b0011010110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010110110000000010) && ({row_reg, col_reg}<22'b0011010110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010110110000101101) && ({row_reg, col_reg}<22'b0011010111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010111000001010111) && ({row_reg, col_reg}<22'b0011010111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010111000010000010) && ({row_reg, col_reg}<22'b0011010111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010111000100000010) && ({row_reg, col_reg}<22'b0011010111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010111000100101101) && ({row_reg, col_reg}<22'b0011010111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010111001101010111) && ({row_reg, col_reg}<22'b0011010111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011010111001110000010) && ({row_reg, col_reg}<22'b0011010111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010111010000000010) && ({row_reg, col_reg}<22'b0011010111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010111010000101101) && ({row_reg, col_reg}<22'b0011010111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010111100001010111) && ({row_reg, col_reg}<22'b0011010111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011010111100010000010) && ({row_reg, col_reg}<22'b0011010111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010111100100000010) && ({row_reg, col_reg}<22'b0011010111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010111100100101101) && ({row_reg, col_reg}<22'b0011010111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011010111101101010111) && ({row_reg, col_reg}<22'b0011010111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011010111101110000010) && ({row_reg, col_reg}<22'b0011010111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011010111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011010111110000000010) && ({row_reg, col_reg}<22'b0011010111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011010111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011010111110000101101) && ({row_reg, col_reg}<22'b0011011000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011000000001010111) && ({row_reg, col_reg}<22'b0011011000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011000000010000010) && ({row_reg, col_reg}<22'b0011011000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011000000100000010) && ({row_reg, col_reg}<22'b0011011000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011000000100101101) && ({row_reg, col_reg}<22'b0011011000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011000001101010111) && ({row_reg, col_reg}<22'b0011011000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011011000001110000010) && ({row_reg, col_reg}<22'b0011011000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011000010000000010) && ({row_reg, col_reg}<22'b0011011000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011000010000101101) && ({row_reg, col_reg}<22'b0011011000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011000100001010111) && ({row_reg, col_reg}<22'b0011011000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011000100010000010) && ({row_reg, col_reg}<22'b0011011000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011000100100000010) && ({row_reg, col_reg}<22'b0011011000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011000100100101101) && ({row_reg, col_reg}<22'b0011011000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011000101101010111) && ({row_reg, col_reg}<22'b0011011000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011011000101110000010) && ({row_reg, col_reg}<22'b0011011000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011000110000000010) && ({row_reg, col_reg}<22'b0011011000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011000110000101101) && ({row_reg, col_reg}<22'b0011011001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011001000001010111) && ({row_reg, col_reg}<22'b0011011001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011001000010000010) && ({row_reg, col_reg}<22'b0011011001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011001000100000010) && ({row_reg, col_reg}<22'b0011011001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011001000100101101) && ({row_reg, col_reg}<22'b0011011001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011001001101010111) && ({row_reg, col_reg}<22'b0011011001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011011001001110000010) && ({row_reg, col_reg}<22'b0011011001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011001010000000010) && ({row_reg, col_reg}<22'b0011011001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011001010000101101) && ({row_reg, col_reg}<22'b0011011001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011001100001010111) && ({row_reg, col_reg}<22'b0011011001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011001100010000010) && ({row_reg, col_reg}<22'b0011011001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011001100100000010) && ({row_reg, col_reg}<22'b0011011001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011001100100101101) && ({row_reg, col_reg}<22'b0011011001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011001101101010111) && ({row_reg, col_reg}<22'b0011011001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011001101110000010) && ({row_reg, col_reg}<22'b0011011001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011001110000000010) && ({row_reg, col_reg}<22'b0011011001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011001110000101101) && ({row_reg, col_reg}<22'b0011011010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011010000001010111) && ({row_reg, col_reg}<22'b0011011010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011011010000010000010) && ({row_reg, col_reg}<22'b0011011010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011010000100000010) && ({row_reg, col_reg}<22'b0011011010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011010000100101101) && ({row_reg, col_reg}<22'b0011011010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011010001101010111) && ({row_reg, col_reg}<22'b0011011010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011010001110000010) && ({row_reg, col_reg}<22'b0011011010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011010010000000010) && ({row_reg, col_reg}<22'b0011011010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011010010000101101) && ({row_reg, col_reg}<22'b0011011010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011010100001010111) && ({row_reg, col_reg}<22'b0011011010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011011010100010000010) && ({row_reg, col_reg}<22'b0011011010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011010100100000010) && ({row_reg, col_reg}<22'b0011011010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011010100100101101) && ({row_reg, col_reg}<22'b0011011010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011010101101010111) && ({row_reg, col_reg}<22'b0011011010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011010101110000010) && ({row_reg, col_reg}<22'b0011011010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011010110000000010) && ({row_reg, col_reg}<22'b0011011010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011010110000101101) && ({row_reg, col_reg}<22'b0011011011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011011000001010111) && ({row_reg, col_reg}<22'b0011011011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011011011000010000010) && ({row_reg, col_reg}<22'b0011011011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011011000100000010) && ({row_reg, col_reg}<22'b0011011011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011011000100101101) && ({row_reg, col_reg}<22'b0011011011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011011001101010111) && ({row_reg, col_reg}<22'b0011011011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011011001110000010) && ({row_reg, col_reg}<22'b0011011011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011011010000000010) && ({row_reg, col_reg}<22'b0011011011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011011010000101101) && ({row_reg, col_reg}<22'b0011011011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011011100001010111) && ({row_reg, col_reg}<22'b0011011011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011011011100010000010) && ({row_reg, col_reg}<22'b0011011011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011011100100000010) && ({row_reg, col_reg}<22'b0011011011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011011100100101101) && ({row_reg, col_reg}<22'b0011011011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011011101101010111) && ({row_reg, col_reg}<22'b0011011011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011011101110000010) && ({row_reg, col_reg}<22'b0011011011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011011110000000010) && ({row_reg, col_reg}<22'b0011011011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011011110000101101) && ({row_reg, col_reg}<22'b0011011100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011100000001010111) && ({row_reg, col_reg}<22'b0011011100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0011011100000010000010) && ({row_reg, col_reg}<22'b0011011100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011100000100000010) && ({row_reg, col_reg}<22'b0011011100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011100000100101101) && ({row_reg, col_reg}<22'b0011011100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011100001101010111) && ({row_reg, col_reg}<22'b0011011100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011100001110000010) && ({row_reg, col_reg}<22'b0011011100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011100010000000010) && ({row_reg, col_reg}<22'b0011011100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011100010000101101) && ({row_reg, col_reg}<22'b0011011100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011100100001010111) && ({row_reg, col_reg}<22'b0011011100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011011100100010000010) && ({row_reg, col_reg}<22'b0011011100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011100100100000010) && ({row_reg, col_reg}<22'b0011011100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011100100100101101) && ({row_reg, col_reg}<22'b0011011100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011100101101010111) && ({row_reg, col_reg}<22'b0011011100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011100101110000010) && ({row_reg, col_reg}<22'b0011011100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011100110000000010) && ({row_reg, col_reg}<22'b0011011100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011100110000101101) && ({row_reg, col_reg}<22'b0011011101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011101000001010111) && ({row_reg, col_reg}<22'b0011011101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0011011101000010000010) && ({row_reg, col_reg}<22'b0011011101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011101000100000010) && ({row_reg, col_reg}<22'b0011011101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011101000100101101) && ({row_reg, col_reg}<22'b0011011101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011101001101010111) && ({row_reg, col_reg}<22'b0011011101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011101001110000010) && ({row_reg, col_reg}<22'b0011011101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011101010000000010) && ({row_reg, col_reg}<22'b0011011101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011101010000101101) && ({row_reg, col_reg}<22'b0011011101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011101100001010111) && ({row_reg, col_reg}<22'b0011011101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011101100010000010) && ({row_reg, col_reg}<22'b0011011101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011101100100000010) && ({row_reg, col_reg}<22'b0011011101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011101100100101101) && ({row_reg, col_reg}<22'b0011011101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011101101101010111) && ({row_reg, col_reg}<22'b0011011101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011101101110000010) && ({row_reg, col_reg}<22'b0011011101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011101110000000010) && ({row_reg, col_reg}<22'b0011011101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011101110000101101) && ({row_reg, col_reg}<22'b0011011110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011110000001010111) && ({row_reg, col_reg}<22'b0011011110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011110000010000010) && ({row_reg, col_reg}<22'b0011011110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011110000100000010) && ({row_reg, col_reg}<22'b0011011110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011110000100101101) && ({row_reg, col_reg}<22'b0011011110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011110001101010111) && ({row_reg, col_reg}<22'b0011011110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011110001110000010) && ({row_reg, col_reg}<22'b0011011110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011110010000000010) && ({row_reg, col_reg}<22'b0011011110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011110010000101101) && ({row_reg, col_reg}<22'b0011011110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011110100001010111) && ({row_reg, col_reg}<22'b0011011110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011110100010000010) && ({row_reg, col_reg}<22'b0011011110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011110100100000010) && ({row_reg, col_reg}<22'b0011011110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011110100100101101) && ({row_reg, col_reg}<22'b0011011110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011110101101010111) && ({row_reg, col_reg}<22'b0011011110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011110101110000010) && ({row_reg, col_reg}<22'b0011011110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011110110000000010) && ({row_reg, col_reg}<22'b0011011110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011110110000101101) && ({row_reg, col_reg}<22'b0011011111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011111000001010111) && ({row_reg, col_reg}<22'b0011011111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011111000010000010) && ({row_reg, col_reg}<22'b0011011111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011111000100000010) && ({row_reg, col_reg}<22'b0011011111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011111000100101101) && ({row_reg, col_reg}<22'b0011011111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011111001101010111) && ({row_reg, col_reg}<22'b0011011111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011111001110000010) && ({row_reg, col_reg}<22'b0011011111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011111010000000010) && ({row_reg, col_reg}<22'b0011011111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011111010000101101) && ({row_reg, col_reg}<22'b0011011111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011111100001010111) && ({row_reg, col_reg}<22'b0011011111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011111100010000010) && ({row_reg, col_reg}<22'b0011011111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011111100100000010) && ({row_reg, col_reg}<22'b0011011111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011111100100101101) && ({row_reg, col_reg}<22'b0011011111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011011111101101010111) && ({row_reg, col_reg}<22'b0011011111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011011111101110000010) && ({row_reg, col_reg}<22'b0011011111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011011111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011011111110000000010) && ({row_reg, col_reg}<22'b0011011111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011011111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011011111110000101101) && ({row_reg, col_reg}<22'b0011100000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100000000001010111) && ({row_reg, col_reg}<22'b0011100000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100000000010000001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=22'b0011100000000010000010) && ({row_reg, col_reg}<22'b0011100000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==22'b0011100000000100000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011100000000100000010) && ({row_reg, col_reg}<22'b0011100000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100000000100101101) && ({row_reg, col_reg}<22'b0011100000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100000001101010111) && ({row_reg, col_reg}<22'b0011100000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100000001110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011100000001110000010) && ({row_reg, col_reg}<22'b0011100000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==22'b0011100000010000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011100000010000000010) && ({row_reg, col_reg}<22'b0011100000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100000010000101101) && ({row_reg, col_reg}<22'b0011100000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100000100001010111) && ({row_reg, col_reg}<22'b0011100000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100000100100101101) && ({row_reg, col_reg}<22'b0011100000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100000101101010111) && ({row_reg, col_reg}<22'b0011100000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100000110000101101) && ({row_reg, col_reg}<22'b0011100001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100001000001010111) && ({row_reg, col_reg}<22'b0011100001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100001000100101101) && ({row_reg, col_reg}<22'b0011100001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100001001101010111) && ({row_reg, col_reg}<22'b0011100001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100001010000101101) && ({row_reg, col_reg}<22'b0011100001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100001100001010111) && ({row_reg, col_reg}<22'b0011100001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100001100100101101) && ({row_reg, col_reg}<22'b0011100001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100001101101010111) && ({row_reg, col_reg}<22'b0011100001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100001110000101101) && ({row_reg, col_reg}<22'b0011100010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100010000001010111) && ({row_reg, col_reg}<22'b0011100010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100010000100101101) && ({row_reg, col_reg}<22'b0011100010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100010001101010111) && ({row_reg, col_reg}<22'b0011100010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100010010000101101) && ({row_reg, col_reg}<22'b0011100010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100010100001010111) && ({row_reg, col_reg}<22'b0011100010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100010100100101101) && ({row_reg, col_reg}<22'b0011100010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100010101101010111) && ({row_reg, col_reg}<22'b0011100010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100010110000101101) && ({row_reg, col_reg}<22'b0011100011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100011000001010111) && ({row_reg, col_reg}<22'b0011100011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100011000100101101) && ({row_reg, col_reg}<22'b0011100011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100011001101010111) && ({row_reg, col_reg}<22'b0011100011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100011010000101101) && ({row_reg, col_reg}<22'b0011100011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100011100001010111) && ({row_reg, col_reg}<22'b0011100011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100011100100101101) && ({row_reg, col_reg}<22'b0011100011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100011101101010111) && ({row_reg, col_reg}<22'b0011100011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100011110000101101) && ({row_reg, col_reg}<22'b0011100100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100100000001010111) && ({row_reg, col_reg}<22'b0011100100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100100000100101101) && ({row_reg, col_reg}<22'b0011100100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100100001101010111) && ({row_reg, col_reg}<22'b0011100100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100100010000101101) && ({row_reg, col_reg}<22'b0011100100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100100100001010111) && ({row_reg, col_reg}<22'b0011100100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100100100100101101) && ({row_reg, col_reg}<22'b0011100100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100100101101010111) && ({row_reg, col_reg}<22'b0011100100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100100110000101101) && ({row_reg, col_reg}<22'b0011100101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100101000001010111) && ({row_reg, col_reg}<22'b0011100101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100101000100101101) && ({row_reg, col_reg}<22'b0011100101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100101001101010111) && ({row_reg, col_reg}<22'b0011100101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100101010000101101) && ({row_reg, col_reg}<22'b0011100101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100101100001010111) && ({row_reg, col_reg}<22'b0011100101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100101100100101101) && ({row_reg, col_reg}<22'b0011100101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100101101101010111) && ({row_reg, col_reg}<22'b0011100101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100101110000101101) && ({row_reg, col_reg}<22'b0011100110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100110000001010111) && ({row_reg, col_reg}<22'b0011100110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100110000100101101) && ({row_reg, col_reg}<22'b0011100110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100110001101010111) && ({row_reg, col_reg}<22'b0011100110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100110010000101101) && ({row_reg, col_reg}<22'b0011100110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100110100001010111) && ({row_reg, col_reg}<22'b0011100110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100110100100101101) && ({row_reg, col_reg}<22'b0011100110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100110101101010111) && ({row_reg, col_reg}<22'b0011100110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100110110000101101) && ({row_reg, col_reg}<22'b0011100111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100111000001010111) && ({row_reg, col_reg}<22'b0011100111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100111000100101101) && ({row_reg, col_reg}<22'b0011100111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100111001101010111) && ({row_reg, col_reg}<22'b0011100111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100111010000101101) && ({row_reg, col_reg}<22'b0011100111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100111100001010111) && ({row_reg, col_reg}<22'b0011100111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011100111100100101101) && ({row_reg, col_reg}<22'b0011100111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011100111101101010111) && ({row_reg, col_reg}<22'b0011100111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011100111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011100111110000101101) && ({row_reg, col_reg}<22'b0011101000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101000000001010111) && ({row_reg, col_reg}<22'b0011101000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011101000000100101101) && ({row_reg, col_reg}<22'b0011101000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101000001101010111) && ({row_reg, col_reg}<22'b0011101000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011101000010000101101) && ({row_reg, col_reg}<22'b0011101000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101000100001010111) && ({row_reg, col_reg}<22'b0011101000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011101000100100101101) && ({row_reg, col_reg}<22'b0011101000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101000101101010111) && ({row_reg, col_reg}<22'b0011101000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011101000110000101101) && ({row_reg, col_reg}<22'b0011101001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101001000001010111) && ({row_reg, col_reg}<22'b0011101001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011101001000100101101) && ({row_reg, col_reg}<22'b0011101001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101001001101010111) && ({row_reg, col_reg}<22'b0011101001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011101001010000101101) && ({row_reg, col_reg}<22'b0011101001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101001100001010111) && ({row_reg, col_reg}<22'b0011101001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011101001100100101101) && ({row_reg, col_reg}<22'b0011101001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101001101101010111) && ({row_reg, col_reg}<22'b0011101001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011101001110000101101) && ({row_reg, col_reg}<22'b0011101010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101010000001010111) && ({row_reg, col_reg}<22'b0011101010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011101010000100101101) && ({row_reg, col_reg}<22'b0011101010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101010001101010111) && ({row_reg, col_reg}<22'b0011101010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011101010010000101101) && ({row_reg, col_reg}<22'b0011101010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101010100001010111) && ({row_reg, col_reg}<22'b0011101010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011101010100100101101) && ({row_reg, col_reg}<22'b0011101010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101010101101010111) && ({row_reg, col_reg}<22'b0011101010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011101010110000101101) && ({row_reg, col_reg}<22'b0011101011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101011000001010111) && ({row_reg, col_reg}<22'b0011101011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011101011000100101101) && ({row_reg, col_reg}<22'b0011101011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101011001101010111) && ({row_reg, col_reg}<22'b0011101011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0011101011010000101101) && ({row_reg, col_reg}<22'b0011101011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101011100001010111) && ({row_reg, col_reg}<22'b0011101011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011101011100100101100) && ({row_reg, col_reg}<22'b0011101011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101011101101010111) && ({row_reg, col_reg}<22'b0011101011110000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011101011110000101100) && ({row_reg, col_reg}<22'b0011101100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101100000001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011101100000001011000) && ({row_reg, col_reg}<22'b0011101100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011101100000100101100) && ({row_reg, col_reg}<22'b0011101100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101100001101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011101100001101011000) && ({row_reg, col_reg}<22'b0011101100010000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011101100010000101100) && ({row_reg, col_reg}<22'b0011101100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101100100001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0011101100100001011000) && ({row_reg, col_reg}<22'b0011101100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011101100100100101100) && ({row_reg, col_reg}<22'b0011101100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101100101101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0011101100101101011000) && ({row_reg, col_reg}<22'b0011101100110000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011101100110000101100) && ({row_reg, col_reg}<22'b0011101101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101101000001010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011101101000001011000) && ({row_reg, col_reg}<22'b0011101101000100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101101000100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011101101000100101100) && ({row_reg, col_reg}<22'b0011101101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101101001101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011101101001101011000) && ({row_reg, col_reg}<22'b0011101101010000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101101010000101011)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=22'b0011101101010000101100) && ({row_reg, col_reg}<22'b0011101101100001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101101100001011000) && ({row_reg, col_reg}<22'b0011101101100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101101100100101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011101101100100101100) && ({row_reg, col_reg}<22'b0011101101101101011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101101101101011000) && ({row_reg, col_reg}<22'b0011101101110000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101101110000101011)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0011101101110000101100) && ({row_reg, col_reg}<22'b0011101110000001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101110000001011000) && ({row_reg, col_reg}<22'b0011101110000100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011101110000100101011) && ({row_reg, col_reg}<22'b0011101110001101011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101110001101011000) && ({row_reg, col_reg}<22'b0011101110010000101011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011101110010000101011) && ({row_reg, col_reg}<22'b0011101110100001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101110100001011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011101110100001011001) && ({row_reg, col_reg}<22'b0011101110100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011101110100100101011) && ({row_reg, col_reg}<22'b0011101110101101011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101110101101011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011101110101101011001) && ({row_reg, col_reg}<22'b0011101110110000101011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011101110110000101011) && ({row_reg, col_reg}<22'b0011101111000001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101111000001011001) && ({row_reg, col_reg}<22'b0011101111000100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101111000100101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011101111000100101011) && ({row_reg, col_reg}<22'b0011101111001101011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011101111001101011001) && ({row_reg, col_reg}<22'b0011101111010000101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011101111010000101010)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0011101111010000101011) && ({row_reg, col_reg}<22'b0011101111100001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101111100001011001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}>=22'b0011101111100001011010) && ({row_reg, col_reg}<22'b0011101111100100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011101111100100101010) && ({row_reg, col_reg}<22'b0011101111101101011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011101111101101011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0011101111101101011010) && ({row_reg, col_reg}<22'b0011101111110000101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011101111110000101010) && ({row_reg, col_reg}<22'b0011110000000001011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110000000001011010) && ({row_reg, col_reg}<22'b0011110000000100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110000000100101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011110000000100101010) && ({row_reg, col_reg}<22'b0011110000001101011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110000001101011010) && ({row_reg, col_reg}<22'b0011110000010000101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110000010000101001)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0011110000010000101010) && ({row_reg, col_reg}<22'b0011110000100001011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110000100001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011110000100001011011) && ({row_reg, col_reg}<22'b0011110000100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011110000100100101001) && ({row_reg, col_reg}<22'b0011110000101101011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110000101101011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011110000101101011011) && ({row_reg, col_reg}<22'b0011110000110000101001)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011110000110000101001) && ({row_reg, col_reg}<22'b0011110001000001011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110001000001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011110001000001011100) && ({row_reg, col_reg}<22'b0011110001000100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011110001000100101000) && ({row_reg, col_reg}<22'b0011110001001101011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110001001101011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011110001001101011100) && ({row_reg, col_reg}<22'b0011110001010000101000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011110001010000101000) && ({row_reg, col_reg}<22'b0011110001100001011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110001100001011100) && ({row_reg, col_reg}<22'b0011110001100100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110001100100100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011110001100100101000) && ({row_reg, col_reg}<22'b0011110001101101011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110001101101011100) && ({row_reg, col_reg}<22'b0011110001110000100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110001110000100111)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0011110001110000101000) && ({row_reg, col_reg}<22'b0011110010000001011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110010000001011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011110010000001011101) && ({row_reg, col_reg}<22'b0011110010000100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110010000100100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011110010000100100111) && ({row_reg, col_reg}<22'b0011110010001101011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110010001101011100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011110010001101011101) && ({row_reg, col_reg}<22'b0011110010010000100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110010010000100110)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0011110010010000100111) && ({row_reg, col_reg}<22'b0011110010100001011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110010100001011110) && ({row_reg, col_reg}<22'b0011110010100100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110010100100100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011110010100100100110) && ({row_reg, col_reg}<22'b0011110010101101011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110010101101011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011110010101101011110) && ({row_reg, col_reg}<22'b0011110010110000100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110010110000100101)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0011110010110000100110) && ({row_reg, col_reg}<22'b0011110011000001011111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110011000001011111) && ({row_reg, col_reg}<22'b0011110011000100100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110011000100100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011110011000100100101) && ({row_reg, col_reg}<22'b0011110011001101011111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110011001101011111) && ({row_reg, col_reg}<22'b0011110011010000100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110011010000100100)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0011110011010000100101) && ({row_reg, col_reg}<22'b0011110011100001100000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110011100001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0011110011100001100001) && ({row_reg, col_reg}<22'b0011110011100100100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0011110011100100100011) && ({row_reg, col_reg}<22'b0011110011101101100000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110011101101100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0011110011101101100001) && ({row_reg, col_reg}<22'b0011110011110000100011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0011110011110000100011) && ({row_reg, col_reg}<22'b0011110100000001100001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110100000001100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011110100000001100010) && ({row_reg, col_reg}<22'b0011110100000100100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110100000100100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011110100000100100010) && ({row_reg, col_reg}<22'b0011110100001101100001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110100001101100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==22'b0011110100001101100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0011110100001101100011) && ({row_reg, col_reg}<22'b0011110100010000100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110100010000100001)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0011110100010000100010) && ({row_reg, col_reg}<22'b0011110100100001100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110100100001100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==22'b0011110100100001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011110100100001100101) && ({row_reg, col_reg}<22'b0011110100100100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110100100100011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0011110100100100100000) && ({row_reg, col_reg}<22'b0011110100101101100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110100101101100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==22'b0011110100101101100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0011110100101101100101) && ({row_reg, col_reg}<22'b0011110100110000011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110100110000011111)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0011110100110000100000) && ({row_reg, col_reg}<22'b0011110101000001100110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110101000001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0011110101000001100111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=22'b0011110101000001101000) && ({row_reg, col_reg}<22'b0011110101000100011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110101000100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==22'b0011110101000100011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0011110101000100011101) && ({row_reg, col_reg}<22'b0011110101001101100110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0011110101001101100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0011110101001101100111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=22'b0011110101001101101000) && ({row_reg, col_reg}<22'b0011110101010000011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0011110101010000011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==22'b0011110101010000011100)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0011110101010000011101) && ({row_reg, col_reg}<22'b0011110101100001101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110101100001101011) && ({row_reg, col_reg}<22'b0011110101100100011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0011110101100100011000) && ({row_reg, col_reg}<22'b0011110101101101101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0011110101101101101011) && ({row_reg, col_reg}<22'b0011110101110000011000)) color_data = 12'b110011001100;
































































































































		if(({row_reg, col_reg}>=22'b0011110101110000011000) && ({row_reg, col_reg}<22'b0100110101100001101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110101100001101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==22'b0100110101100001101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0100110101100001101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100001101100) && ({row_reg, col_reg}<22'b0100110101100001110001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100001110001) && ({row_reg, col_reg}<22'b0100110101100001111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100001111110) && ({row_reg, col_reg}<22'b0100110101100010000101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100010000101) && ({row_reg, col_reg}<22'b0100110101100010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100010010010) && ({row_reg, col_reg}<22'b0100110101100010011001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100010011001) && ({row_reg, col_reg}<22'b0100110101100010100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100010100110) && ({row_reg, col_reg}<22'b0100110101100010101101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100010101101) && ({row_reg, col_reg}<22'b0100110101100010111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100010111010) && ({row_reg, col_reg}<22'b0100110101100011000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100011000001) && ({row_reg, col_reg}<22'b0100110101100011001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100011001110) && ({row_reg, col_reg}<22'b0100110101100011010101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100011010101) && ({row_reg, col_reg}<22'b0100110101100011100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100011100010) && ({row_reg, col_reg}<22'b0100110101100011101001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100011101001) && ({row_reg, col_reg}<22'b0100110101100011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100011110110) && ({row_reg, col_reg}<22'b0100110101100011111101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100011111101) && ({row_reg, col_reg}<22'b0100110101100100001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101100100001010) && ({row_reg, col_reg}<22'b0100110101100100010001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101100100010001) && ({row_reg, col_reg}<22'b0100110101100100011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b0100110101100100011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0100110101100100011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0100110101100100011011) && ({row_reg, col_reg}<22'b0100110101101101101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110101101101101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==22'b0100110101101101101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0100110101101101101011) && ({row_reg, col_reg}<22'b0100110101101101110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101101101110110) && ({row_reg, col_reg}<22'b0100110101101101111101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101101101111101) && ({row_reg, col_reg}<22'b0100110101101110001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101101110001010) && ({row_reg, col_reg}<22'b0100110101101110010001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101101110010001) && ({row_reg, col_reg}<22'b0100110101101110011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101101110011110) && ({row_reg, col_reg}<22'b0100110101101110100101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101101110100101) && ({row_reg, col_reg}<22'b0100110101101110110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101101110110010) && ({row_reg, col_reg}<22'b0100110101101110111001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101101110111001) && ({row_reg, col_reg}<22'b0100110101101111000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101101111000110) && ({row_reg, col_reg}<22'b0100110101101111001101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101101111001101) && ({row_reg, col_reg}<22'b0100110101101111011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101101111011010) && ({row_reg, col_reg}<22'b0100110101101111100001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101101111100001) && ({row_reg, col_reg}<22'b0100110101101111101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101101111101110) && ({row_reg, col_reg}<22'b0100110101101111110101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101101111110101) && ({row_reg, col_reg}<22'b0100110101110000000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101110000000010) && ({row_reg, col_reg}<22'b0100110101110000001001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0100110101110000001001) && ({row_reg, col_reg}<22'b0100110101110000010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110101110000010110) && ({row_reg, col_reg}<22'b0100110101110000011000)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==22'b0100110101110000011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b0100110101110000011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0100110101110000011010)) color_data = 12'b101110111100;

		if(({row_reg, col_reg}>=22'b0100110101110000011011) && ({row_reg, col_reg}<22'b0100110110000001100101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110110000001100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0100110110000001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0100110110000001100111) && ({row_reg, col_reg}<22'b0100110110000100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110110000100011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110110000100011110) && ({row_reg, col_reg}<22'b0100110110001101100101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110110001101100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b0100110110001101100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0100110110001101100111) && ({row_reg, col_reg}<22'b0100110110010000011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110110010000011101)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0100110110010000011110) && ({row_reg, col_reg}<22'b0100110110100001100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110110100001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100110110100001100100) && ({row_reg, col_reg}<22'b0100110110100100011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110110100100011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==22'b0100110110100100100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0100110110100100100001) && ({row_reg, col_reg}<22'b0100110110101101100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110110101101100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100110110101101100100) && ({row_reg, col_reg}<22'b0100110110110000011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110110110000011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==22'b0100110110110000100000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=22'b0100110110110000100001) && ({row_reg, col_reg}<22'b0100110111000001100001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110111000001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100110111000001100010) && ({row_reg, col_reg}<22'b0100110111000100100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110111000100100001)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0100110111000100100010) && ({row_reg, col_reg}<22'b0100110111001101100001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110111001101100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100110111001101100010) && ({row_reg, col_reg}<22'b0100110111010000100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110111010000100001)) color_data = 12'b011001100111;

		if(({row_reg, col_reg}>=22'b0100110111010000100010) && ({row_reg, col_reg}<22'b0100110111100001011111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110111100001011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0100110111100001100000) && ({row_reg, col_reg}<22'b0100110111100100100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110111100100100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100110111100100100100) && ({row_reg, col_reg}<22'b0100110111101101011111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100110111101101011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0100110111101101100000) && ({row_reg, col_reg}<22'b0100110111110000100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100110111110000100011)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b0100110111110000100100) && ({row_reg, col_reg}<22'b0100111000000001011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111000000001011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0100111000000001011111) && ({row_reg, col_reg}<22'b0100111000000100100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111000000100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0100111000000100100101) && ({row_reg, col_reg}<22'b0100111000001101011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111000001101011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0100111000001101011111) && ({row_reg, col_reg}<22'b0100111000010000100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111000010000100100)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=22'b0100111000010000100101) && ({row_reg, col_reg}<22'b0100111000100001011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111000100001011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100111000100001011110) && ({row_reg, col_reg}<22'b0100111000100100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111000100100100101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=22'b0100111000100100100110) && ({row_reg, col_reg}<22'b0100111000101101011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111000101101011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100111000101101011110) && ({row_reg, col_reg}<22'b0100111000110000100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111000110000100101)) color_data = 12'b011001100111;

		if(({row_reg, col_reg}>=22'b0100111000110000100110) && ({row_reg, col_reg}<22'b0100111001000001011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111001000001011100)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=22'b0100111001000001011101) && ({row_reg, col_reg}<22'b0100111001000100100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111001000100100110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=22'b0100111001000100100111) && ({row_reg, col_reg}<22'b0100111001001101011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111001001101011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100111001001101011101) && ({row_reg, col_reg}<22'b0100111001010000100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111001010000100110)) color_data = 12'b011001100111;

		if(({row_reg, col_reg}>=22'b0100111001010000100111) && ({row_reg, col_reg}<22'b0100111001100001011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111001100001011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0100111001100001011100) && ({row_reg, col_reg}<22'b0100111001100100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111001100100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100111001100100101000) && ({row_reg, col_reg}<22'b0100111001101101011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111001101101011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0100111001101101011100) && ({row_reg, col_reg}<22'b0100111001110000100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111001110000100111)) color_data = 12'b011110001000;

		if(({row_reg, col_reg}>=22'b0100111001110000101000) && ({row_reg, col_reg}<22'b0100111010000001011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111010000001011011) && ({row_reg, col_reg}<22'b0100111010000100101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111010000100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0100111010000100101001) && ({row_reg, col_reg}<22'b0100111010001101011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111010001101011011) && ({row_reg, col_reg}<22'b0100111010010000101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111010010000101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b0100111010010000101001) && ({row_reg, col_reg}<22'b0100111010100001011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111010100001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0100111010100001011011) && ({row_reg, col_reg}<22'b0100111010100100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0100111010100100101001) && ({row_reg, col_reg}<22'b0100111010101101011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111010101101011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0100111010101101011011) && ({row_reg, col_reg}<22'b0100111010110000101001)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0100111010110000101001) && ({row_reg, col_reg}<22'b0100111011000001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111011000001011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0100111011000001011010) && ({row_reg, col_reg}<22'b0100111011000100101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111011000100101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100111011000100101010) && ({row_reg, col_reg}<22'b0100111011001101011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111011001101011001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0100111011001101011010) && ({row_reg, col_reg}<22'b0100111011010000101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111011010000101001)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=22'b0100111011010000101010) && ({row_reg, col_reg}<22'b0100111011100001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111011100001011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0100111011100001011010) && ({row_reg, col_reg}<22'b0100111011100100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0100111011100100101010) && ({row_reg, col_reg}<22'b0100111011101101011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111011101101011001) && ({row_reg, col_reg}<22'b0100111011110000101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0100111011110000101010) && ({row_reg, col_reg}<22'b0100111100000001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111100000001011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0100111100000001011001) && ({row_reg, col_reg}<22'b0100111100000100101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111100000100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100111100000100101011) && ({row_reg, col_reg}<22'b0100111100001101011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111100001101011000)) color_data = 12'b101110111100;
		if(({row_reg, col_reg}>=22'b0100111100001101011001) && ({row_reg, col_reg}<22'b0100111100010000101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111100010000101010)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=22'b0100111100010000101011) && ({row_reg, col_reg}<22'b0100111100100001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111100100001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100111100100001011001) && ({row_reg, col_reg}<22'b0100111100100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0100111100100100101011) && ({row_reg, col_reg}<22'b0100111100101101011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111100101101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100111100101101011001) && ({row_reg, col_reg}<22'b0100111100110000101011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0100111100110000101011) && ({row_reg, col_reg}<22'b0100111101000001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111101000001011000) && ({row_reg, col_reg}<22'b0100111101000100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111101000100101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0100111101000100101100) && ({row_reg, col_reg}<22'b0100111101001101011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111101001101011000) && ({row_reg, col_reg}<22'b0100111101010000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111101010000101011)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=22'b0100111101010000101100) && ({row_reg, col_reg}<22'b0100111101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111101100001010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0100111101100001011000) && ({row_reg, col_reg}<22'b0100111101100100101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111101100100101011)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0100111101100100101100) && ({row_reg, col_reg}<22'b0100111101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111101101101010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0100111101101101011000) && ({row_reg, col_reg}<22'b0100111101110000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0100111101110000101011)) color_data = 12'b100010011001;

		if(({row_reg, col_reg}>=22'b0100111101110000101100) && ({row_reg, col_reg}<22'b0100111110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111110000001010111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=22'b0100111110000001011000) && ({row_reg, col_reg}<22'b0100111110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0100111110000100101100) && ({row_reg, col_reg}<22'b0100111110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111110001101010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0100111110001101011000) && ({row_reg, col_reg}<22'b0100111110010000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0100111110010000101100) && ({row_reg, col_reg}<22'b0100111110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111110100001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100111110100001011000) && ({row_reg, col_reg}<22'b0100111110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0100111110100100101100) && ({row_reg, col_reg}<22'b0100111110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111110101101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0100111110101101011000) && ({row_reg, col_reg}<22'b0100111110110000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0100111110110000101100) && ({row_reg, col_reg}<22'b0100111111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111111000001010111) && ({row_reg, col_reg}<22'b0100111111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0100111111000100101100) && ({row_reg, col_reg}<22'b0100111111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0100111111001101010111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0100111111001101011000) && ({row_reg, col_reg}<22'b0100111111010000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0100111111010000101100) && ({row_reg, col_reg}<22'b0100111111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111111100001010111) && ({row_reg, col_reg}<22'b0100111111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0100111111100100101100) && ({row_reg, col_reg}<22'b0100111111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0100111111101101010111) && ({row_reg, col_reg}<22'b0100111111110000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b0100111111110000101100) && ({row_reg, col_reg}<22'b0101000000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000000000001010111) && ({row_reg, col_reg}<22'b0101000000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000000000100101101) && ({row_reg, col_reg}<22'b0101000000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000000001101010111) && ({row_reg, col_reg}<22'b0101000000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000000010000101101) && ({row_reg, col_reg}<22'b0101000000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000000100001010111) && ({row_reg, col_reg}<22'b0101000000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000000100100101101) && ({row_reg, col_reg}<22'b0101000000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000000101101010111) && ({row_reg, col_reg}<22'b0101000000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000000110000101101) && ({row_reg, col_reg}<22'b0101000001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000001000001010111) && ({row_reg, col_reg}<22'b0101000001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000001000100101101) && ({row_reg, col_reg}<22'b0101000001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000001001101010111) && ({row_reg, col_reg}<22'b0101000001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000001010000101101) && ({row_reg, col_reg}<22'b0101000001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000001100001010111) && ({row_reg, col_reg}<22'b0101000001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000001100100101101) && ({row_reg, col_reg}<22'b0101000001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000001101101010111) && ({row_reg, col_reg}<22'b0101000001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000001110000101101) && ({row_reg, col_reg}<22'b0101000010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000010000001010111) && ({row_reg, col_reg}<22'b0101000010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000010000100101101) && ({row_reg, col_reg}<22'b0101000010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000010001101010111) && ({row_reg, col_reg}<22'b0101000010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000010010000101101) && ({row_reg, col_reg}<22'b0101000010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000010100001010111) && ({row_reg, col_reg}<22'b0101000010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000010100100101101) && ({row_reg, col_reg}<22'b0101000010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000010101101010111) && ({row_reg, col_reg}<22'b0101000010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000010110000101101) && ({row_reg, col_reg}<22'b0101000011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000011000001010111) && ({row_reg, col_reg}<22'b0101000011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000011000100101101) && ({row_reg, col_reg}<22'b0101000011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000011001101010111) && ({row_reg, col_reg}<22'b0101000011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000011010000101101) && ({row_reg, col_reg}<22'b0101000011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000011100001010111) && ({row_reg, col_reg}<22'b0101000011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000011100100101101) && ({row_reg, col_reg}<22'b0101000011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000011101101010111) && ({row_reg, col_reg}<22'b0101000011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000011110000101101) && ({row_reg, col_reg}<22'b0101000100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000100000001010111) && ({row_reg, col_reg}<22'b0101000100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000100000100101101) && ({row_reg, col_reg}<22'b0101000100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000100001101010111) && ({row_reg, col_reg}<22'b0101000100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000100010000101101) && ({row_reg, col_reg}<22'b0101000100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000100100001010111) && ({row_reg, col_reg}<22'b0101000100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000100100100101101) && ({row_reg, col_reg}<22'b0101000100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000100101101010111) && ({row_reg, col_reg}<22'b0101000100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000100110000101101) && ({row_reg, col_reg}<22'b0101000101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000101000001010111) && ({row_reg, col_reg}<22'b0101000101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000101000100101101) && ({row_reg, col_reg}<22'b0101000101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000101001101010111) && ({row_reg, col_reg}<22'b0101000101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000101010000101101) && ({row_reg, col_reg}<22'b0101000101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000101100001010111) && ({row_reg, col_reg}<22'b0101000101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000101100100101101) && ({row_reg, col_reg}<22'b0101000101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000101101101010111) && ({row_reg, col_reg}<22'b0101000101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000101110000101101) && ({row_reg, col_reg}<22'b0101000110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000110000001010111) && ({row_reg, col_reg}<22'b0101000110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000110000100101101) && ({row_reg, col_reg}<22'b0101000110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000110001101010111) && ({row_reg, col_reg}<22'b0101000110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000110010000101101) && ({row_reg, col_reg}<22'b0101000110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000110100001010111) && ({row_reg, col_reg}<22'b0101000110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000110100100101101) && ({row_reg, col_reg}<22'b0101000110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000110101101010111) && ({row_reg, col_reg}<22'b0101000110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000110110000101101) && ({row_reg, col_reg}<22'b0101000111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000111000001010111) && ({row_reg, col_reg}<22'b0101000111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000111000100101101) && ({row_reg, col_reg}<22'b0101000111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000111001101010111) && ({row_reg, col_reg}<22'b0101000111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000111010000101101) && ({row_reg, col_reg}<22'b0101000111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000111100001010111) && ({row_reg, col_reg}<22'b0101000111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101000111100100101101) && ({row_reg, col_reg}<22'b0101000111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101000111101101010111) && ({row_reg, col_reg}<22'b0101000111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101000111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101000111110000101101) && ({row_reg, col_reg}<22'b0101001000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001000000001010111) && ({row_reg, col_reg}<22'b0101001000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001000000100101101) && ({row_reg, col_reg}<22'b0101001000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001000001101010111) && ({row_reg, col_reg}<22'b0101001000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001000010000101101) && ({row_reg, col_reg}<22'b0101001000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001000100001010111) && ({row_reg, col_reg}<22'b0101001000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001000100100101101) && ({row_reg, col_reg}<22'b0101001000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001000101101010111) && ({row_reg, col_reg}<22'b0101001000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001000110000101101) && ({row_reg, col_reg}<22'b0101001001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001001000001010111) && ({row_reg, col_reg}<22'b0101001001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001001000100101101) && ({row_reg, col_reg}<22'b0101001001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001001001101010111) && ({row_reg, col_reg}<22'b0101001001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001001010000101101) && ({row_reg, col_reg}<22'b0101001001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001001100001010111) && ({row_reg, col_reg}<22'b0101001001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001001100100101101) && ({row_reg, col_reg}<22'b0101001001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001001101101010111) && ({row_reg, col_reg}<22'b0101001001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001001110000101101) && ({row_reg, col_reg}<22'b0101001010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001010000001010111) && ({row_reg, col_reg}<22'b0101001010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001010000100101101) && ({row_reg, col_reg}<22'b0101001010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001010001101010111) && ({row_reg, col_reg}<22'b0101001010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001010010000101101) && ({row_reg, col_reg}<22'b0101001010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001010100001010111) && ({row_reg, col_reg}<22'b0101001010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001010100100101101) && ({row_reg, col_reg}<22'b0101001010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001010101101010111) && ({row_reg, col_reg}<22'b0101001010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001010110000101101) && ({row_reg, col_reg}<22'b0101001011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001011000001010111) && ({row_reg, col_reg}<22'b0101001011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101001011000010000010) && ({row_reg, col_reg}<22'b0101001011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001011000100000010) && ({row_reg, col_reg}<22'b0101001011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001011000100101101) && ({row_reg, col_reg}<22'b0101001011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001011001101010111) && ({row_reg, col_reg}<22'b0101001011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001011001110000010) && ({row_reg, col_reg}<22'b0101001011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001011010000000010) && ({row_reg, col_reg}<22'b0101001011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001011010000101101) && ({row_reg, col_reg}<22'b0101001011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001011100001010111) && ({row_reg, col_reg}<22'b0101001011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001011100010000010) && ({row_reg, col_reg}<22'b0101001011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001011100100000010) && ({row_reg, col_reg}<22'b0101001011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001011100100101101) && ({row_reg, col_reg}<22'b0101001011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001011101101010111) && ({row_reg, col_reg}<22'b0101001011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001011101110000010) && ({row_reg, col_reg}<22'b0101001011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001011110000000010) && ({row_reg, col_reg}<22'b0101001011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001011110000101101) && ({row_reg, col_reg}<22'b0101001100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001100000001010111) && ({row_reg, col_reg}<22'b0101001100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001100000010000010) && ({row_reg, col_reg}<22'b0101001100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001100000100000010) && ({row_reg, col_reg}<22'b0101001100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001100000100101101) && ({row_reg, col_reg}<22'b0101001100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001100001101010111) && ({row_reg, col_reg}<22'b0101001100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001100001110000010) && ({row_reg, col_reg}<22'b0101001100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001100010000000010) && ({row_reg, col_reg}<22'b0101001100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001100010000101101) && ({row_reg, col_reg}<22'b0101001100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001100100001010111) && ({row_reg, col_reg}<22'b0101001100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001100100010000010) && ({row_reg, col_reg}<22'b0101001100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001100100100000010) && ({row_reg, col_reg}<22'b0101001100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001100100100101101) && ({row_reg, col_reg}<22'b0101001100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001100101101010111) && ({row_reg, col_reg}<22'b0101001100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001100101110000010) && ({row_reg, col_reg}<22'b0101001100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001100110000000010) && ({row_reg, col_reg}<22'b0101001100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001100110000101101) && ({row_reg, col_reg}<22'b0101001101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001101000001010111) && ({row_reg, col_reg}<22'b0101001101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001101000010000010) && ({row_reg, col_reg}<22'b0101001101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001101000100000010) && ({row_reg, col_reg}<22'b0101001101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001101000100101101) && ({row_reg, col_reg}<22'b0101001101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001101001101010111) && ({row_reg, col_reg}<22'b0101001101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001101001110000010) && ({row_reg, col_reg}<22'b0101001101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001101010000000010) && ({row_reg, col_reg}<22'b0101001101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001101010000101101) && ({row_reg, col_reg}<22'b0101001101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001101100001010111) && ({row_reg, col_reg}<22'b0101001101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001101100010000010) && ({row_reg, col_reg}<22'b0101001101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001101100100000010) && ({row_reg, col_reg}<22'b0101001101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001101100100101101) && ({row_reg, col_reg}<22'b0101001101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001101101101010111) && ({row_reg, col_reg}<22'b0101001101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001101101110000010) && ({row_reg, col_reg}<22'b0101001101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001101110000000010) && ({row_reg, col_reg}<22'b0101001101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001101110000101101) && ({row_reg, col_reg}<22'b0101001110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001110000001010111) && ({row_reg, col_reg}<22'b0101001110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001110000010000010) && ({row_reg, col_reg}<22'b0101001110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001110000100000010) && ({row_reg, col_reg}<22'b0101001110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001110000100101101) && ({row_reg, col_reg}<22'b0101001110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001110001101010111) && ({row_reg, col_reg}<22'b0101001110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101001110001110000010) && ({row_reg, col_reg}<22'b0101001110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001110010000000010) && ({row_reg, col_reg}<22'b0101001110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001110010000101101) && ({row_reg, col_reg}<22'b0101001110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001110100001010111) && ({row_reg, col_reg}<22'b0101001110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001110100010000010) && ({row_reg, col_reg}<22'b0101001110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001110100100000010) && ({row_reg, col_reg}<22'b0101001110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001110100100101101) && ({row_reg, col_reg}<22'b0101001110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001110101101010111) && ({row_reg, col_reg}<22'b0101001110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101001110101110000010) && ({row_reg, col_reg}<22'b0101001110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001110110000000010) && ({row_reg, col_reg}<22'b0101001110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001110110000101101) && ({row_reg, col_reg}<22'b0101001111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001111000001010111) && ({row_reg, col_reg}<22'b0101001111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001111000010000010) && ({row_reg, col_reg}<22'b0101001111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001111000100000010) && ({row_reg, col_reg}<22'b0101001111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001111000100101101) && ({row_reg, col_reg}<22'b0101001111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001111001101010111) && ({row_reg, col_reg}<22'b0101001111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101001111001110000010) && ({row_reg, col_reg}<22'b0101001111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001111010000000010) && ({row_reg, col_reg}<22'b0101001111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001111010000101101) && ({row_reg, col_reg}<22'b0101001111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001111100001010111) && ({row_reg, col_reg}<22'b0101001111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101001111100010000010) && ({row_reg, col_reg}<22'b0101001111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001111100100000010) && ({row_reg, col_reg}<22'b0101001111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001111100100101101) && ({row_reg, col_reg}<22'b0101001111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101001111101101010111) && ({row_reg, col_reg}<22'b0101001111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101001111101110000010) && ({row_reg, col_reg}<22'b0101001111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101001111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101001111110000000010) && ({row_reg, col_reg}<22'b0101001111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101001111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101001111110000101101) && ({row_reg, col_reg}<22'b0101010000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010000000001010111) && ({row_reg, col_reg}<22'b0101010000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010000000010000010) && ({row_reg, col_reg}<22'b0101010000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010000000100000010) && ({row_reg, col_reg}<22'b0101010000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010000000100101101) && ({row_reg, col_reg}<22'b0101010000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010000001101010111) && ({row_reg, col_reg}<22'b0101010000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101010000001110000010) && ({row_reg, col_reg}<22'b0101010000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010000010000000010) && ({row_reg, col_reg}<22'b0101010000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010000010000101101) && ({row_reg, col_reg}<22'b0101010000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010000100001010111) && ({row_reg, col_reg}<22'b0101010000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010000100010000010) && ({row_reg, col_reg}<22'b0101010000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010000100100000010) && ({row_reg, col_reg}<22'b0101010000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010000100100101101) && ({row_reg, col_reg}<22'b0101010000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010000101101010111) && ({row_reg, col_reg}<22'b0101010000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101010000101110000010) && ({row_reg, col_reg}<22'b0101010000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010000110000000010) && ({row_reg, col_reg}<22'b0101010000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010000110000101101) && ({row_reg, col_reg}<22'b0101010001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010001000001010111) && ({row_reg, col_reg}<22'b0101010001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010001000010000010) && ({row_reg, col_reg}<22'b0101010001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010001000100000010) && ({row_reg, col_reg}<22'b0101010001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010001000100101101) && ({row_reg, col_reg}<22'b0101010001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010001001101010111) && ({row_reg, col_reg}<22'b0101010001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101010001001110000010) && ({row_reg, col_reg}<22'b0101010001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010001010000000010) && ({row_reg, col_reg}<22'b0101010001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010001010000101101) && ({row_reg, col_reg}<22'b0101010001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010001100001010111) && ({row_reg, col_reg}<22'b0101010001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010001100010000010) && ({row_reg, col_reg}<22'b0101010001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010001100100000010) && ({row_reg, col_reg}<22'b0101010001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010001100100101101) && ({row_reg, col_reg}<22'b0101010001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010001101101010111) && ({row_reg, col_reg}<22'b0101010001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010001101110000010) && ({row_reg, col_reg}<22'b0101010001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010001110000000010) && ({row_reg, col_reg}<22'b0101010001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010001110000101101) && ({row_reg, col_reg}<22'b0101010010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010010000001010111) && ({row_reg, col_reg}<22'b0101010010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101010010000010000010) && ({row_reg, col_reg}<22'b0101010010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010010000100000010) && ({row_reg, col_reg}<22'b0101010010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010010000100101101) && ({row_reg, col_reg}<22'b0101010010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010010001101010111) && ({row_reg, col_reg}<22'b0101010010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010010001110000010) && ({row_reg, col_reg}<22'b0101010010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010010010000000010) && ({row_reg, col_reg}<22'b0101010010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010010010000101101) && ({row_reg, col_reg}<22'b0101010010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010010100001010111) && ({row_reg, col_reg}<22'b0101010010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101010010100010000010) && ({row_reg, col_reg}<22'b0101010010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010010100100000010) && ({row_reg, col_reg}<22'b0101010010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010010100100101101) && ({row_reg, col_reg}<22'b0101010010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010010101101010111) && ({row_reg, col_reg}<22'b0101010010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010010101110000010) && ({row_reg, col_reg}<22'b0101010010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010010110000000010) && ({row_reg, col_reg}<22'b0101010010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010010110000101101) && ({row_reg, col_reg}<22'b0101010011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010011000001010111) && ({row_reg, col_reg}<22'b0101010011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101010011000010000010) && ({row_reg, col_reg}<22'b0101010011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010011000100000010) && ({row_reg, col_reg}<22'b0101010011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010011000100101101) && ({row_reg, col_reg}<22'b0101010011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010011001101010111) && ({row_reg, col_reg}<22'b0101010011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010011001110000010) && ({row_reg, col_reg}<22'b0101010011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010011010000000010) && ({row_reg, col_reg}<22'b0101010011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010011010000101101) && ({row_reg, col_reg}<22'b0101010011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010011100001010111) && ({row_reg, col_reg}<22'b0101010011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101010011100010000010) && ({row_reg, col_reg}<22'b0101010011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010011100100000010) && ({row_reg, col_reg}<22'b0101010011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010011100100101101) && ({row_reg, col_reg}<22'b0101010011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010011101101010111) && ({row_reg, col_reg}<22'b0101010011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010011101110000010) && ({row_reg, col_reg}<22'b0101010011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010011110000000010) && ({row_reg, col_reg}<22'b0101010011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010011110000101101) && ({row_reg, col_reg}<22'b0101010100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010100000001010111) && ({row_reg, col_reg}<22'b0101010100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101010100000010000010) && ({row_reg, col_reg}<22'b0101010100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010100000100000010) && ({row_reg, col_reg}<22'b0101010100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010100000100101101) && ({row_reg, col_reg}<22'b0101010100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010100001101010111) && ({row_reg, col_reg}<22'b0101010100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010100001110000010) && ({row_reg, col_reg}<22'b0101010100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010100010000000010) && ({row_reg, col_reg}<22'b0101010100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010100010000101101) && ({row_reg, col_reg}<22'b0101010100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010100100001010111) && ({row_reg, col_reg}<22'b0101010100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101010100100010000010) && ({row_reg, col_reg}<22'b0101010100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010100100100000010) && ({row_reg, col_reg}<22'b0101010100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010100100100101101) && ({row_reg, col_reg}<22'b0101010100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010100101101010111) && ({row_reg, col_reg}<22'b0101010100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010100101110000010) && ({row_reg, col_reg}<22'b0101010100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010100110000000010) && ({row_reg, col_reg}<22'b0101010100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010100110000101101) && ({row_reg, col_reg}<22'b0101010101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010101000001010111) && ({row_reg, col_reg}<22'b0101010101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101010101000010000010) && ({row_reg, col_reg}<22'b0101010101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010101000100000010) && ({row_reg, col_reg}<22'b0101010101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010101000100101101) && ({row_reg, col_reg}<22'b0101010101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010101001101010111) && ({row_reg, col_reg}<22'b0101010101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010101001110000010) && ({row_reg, col_reg}<22'b0101010101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010101010000000010) && ({row_reg, col_reg}<22'b0101010101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010101010000101101) && ({row_reg, col_reg}<22'b0101010101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010101100001010111) && ({row_reg, col_reg}<22'b0101010101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010101100010000010) && ({row_reg, col_reg}<22'b0101010101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010101100100000010) && ({row_reg, col_reg}<22'b0101010101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010101100100101101) && ({row_reg, col_reg}<22'b0101010101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010101101101010111) && ({row_reg, col_reg}<22'b0101010101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010101101110000010) && ({row_reg, col_reg}<22'b0101010101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010101110000000010) && ({row_reg, col_reg}<22'b0101010101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010101110000101101) && ({row_reg, col_reg}<22'b0101010110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010110000001010111) && ({row_reg, col_reg}<22'b0101010110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010110000010000010) && ({row_reg, col_reg}<22'b0101010110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010110000100000010) && ({row_reg, col_reg}<22'b0101010110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010110000100101101) && ({row_reg, col_reg}<22'b0101010110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010110001101010111) && ({row_reg, col_reg}<22'b0101010110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010110001110000010) && ({row_reg, col_reg}<22'b0101010110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010110010000000010) && ({row_reg, col_reg}<22'b0101010110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010110010000101101) && ({row_reg, col_reg}<22'b0101010110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010110100001010111) && ({row_reg, col_reg}<22'b0101010110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010110100010000010) && ({row_reg, col_reg}<22'b0101010110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010110100100000010) && ({row_reg, col_reg}<22'b0101010110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010110100100101101) && ({row_reg, col_reg}<22'b0101010110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010110101101010111) && ({row_reg, col_reg}<22'b0101010110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010110101110000010) && ({row_reg, col_reg}<22'b0101010110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010110110000000010) && ({row_reg, col_reg}<22'b0101010110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010110110000101101) && ({row_reg, col_reg}<22'b0101010111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010111000001010111) && ({row_reg, col_reg}<22'b0101010111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010111000010000010) && ({row_reg, col_reg}<22'b0101010111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010111000100000010) && ({row_reg, col_reg}<22'b0101010111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010111000100101101) && ({row_reg, col_reg}<22'b0101010111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010111001101010111) && ({row_reg, col_reg}<22'b0101010111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010111001110000010) && ({row_reg, col_reg}<22'b0101010111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010111010000000010) && ({row_reg, col_reg}<22'b0101010111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010111010000101101) && ({row_reg, col_reg}<22'b0101010111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010111100001010111) && ({row_reg, col_reg}<22'b0101010111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010111100010000010) && ({row_reg, col_reg}<22'b0101010111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010111100100000010) && ({row_reg, col_reg}<22'b0101010111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010111100100101101) && ({row_reg, col_reg}<22'b0101010111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101010111101101010111) && ({row_reg, col_reg}<22'b0101010111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101010111101110000010) && ({row_reg, col_reg}<22'b0101010111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101010111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101010111110000000010) && ({row_reg, col_reg}<22'b0101010111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101010111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101010111110000101101) && ({row_reg, col_reg}<22'b0101011000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011000000001010111) && ({row_reg, col_reg}<22'b0101011000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011000000010000010) && ({row_reg, col_reg}<22'b0101011000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011000000100000010) && ({row_reg, col_reg}<22'b0101011000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011000000100101101) && ({row_reg, col_reg}<22'b0101011000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011000001101010111) && ({row_reg, col_reg}<22'b0101011000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011000001110000010) && ({row_reg, col_reg}<22'b0101011000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011000010000000010) && ({row_reg, col_reg}<22'b0101011000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011000010000101101) && ({row_reg, col_reg}<22'b0101011000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011000100001010111) && ({row_reg, col_reg}<22'b0101011000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011000100010000010) && ({row_reg, col_reg}<22'b0101011000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011000100100000010) && ({row_reg, col_reg}<22'b0101011000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011000100100101101) && ({row_reg, col_reg}<22'b0101011000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011000101101010111) && ({row_reg, col_reg}<22'b0101011000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011000101110000010) && ({row_reg, col_reg}<22'b0101011000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011000110000000010) && ({row_reg, col_reg}<22'b0101011000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011000110000101101) && ({row_reg, col_reg}<22'b0101011001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011001000001010111) && ({row_reg, col_reg}<22'b0101011001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011001000010000010) && ({row_reg, col_reg}<22'b0101011001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011001000100000010) && ({row_reg, col_reg}<22'b0101011001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011001000100101101) && ({row_reg, col_reg}<22'b0101011001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011001001101010111) && ({row_reg, col_reg}<22'b0101011001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101011001001110000010) && ({row_reg, col_reg}<22'b0101011001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011001010000000010) && ({row_reg, col_reg}<22'b0101011001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011001010000101101) && ({row_reg, col_reg}<22'b0101011001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011001100001010111) && ({row_reg, col_reg}<22'b0101011001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011001100010000010) && ({row_reg, col_reg}<22'b0101011001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011001100100000010) && ({row_reg, col_reg}<22'b0101011001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011001100100101101) && ({row_reg, col_reg}<22'b0101011001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011001101101010111) && ({row_reg, col_reg}<22'b0101011001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101011001101110000010) && ({row_reg, col_reg}<22'b0101011001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011001110000000010) && ({row_reg, col_reg}<22'b0101011001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011001110000101101) && ({row_reg, col_reg}<22'b0101011010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011010000001010111) && ({row_reg, col_reg}<22'b0101011010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011010000010000010) && ({row_reg, col_reg}<22'b0101011010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011010000100000010) && ({row_reg, col_reg}<22'b0101011010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011010000100101101) && ({row_reg, col_reg}<22'b0101011010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011010001101010111) && ({row_reg, col_reg}<22'b0101011010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101011010001110000010) && ({row_reg, col_reg}<22'b0101011010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011010010000000010) && ({row_reg, col_reg}<22'b0101011010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011010010000101101) && ({row_reg, col_reg}<22'b0101011010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011010100001010111) && ({row_reg, col_reg}<22'b0101011010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011010100010000010) && ({row_reg, col_reg}<22'b0101011010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011010100100000010) && ({row_reg, col_reg}<22'b0101011010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011010100100101101) && ({row_reg, col_reg}<22'b0101011010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011010101101010111) && ({row_reg, col_reg}<22'b0101011010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011010101110000010) && ({row_reg, col_reg}<22'b0101011010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011010110000000010) && ({row_reg, col_reg}<22'b0101011010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011010110000101101) && ({row_reg, col_reg}<22'b0101011011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011011000001010111) && ({row_reg, col_reg}<22'b0101011011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011011000010000010) && ({row_reg, col_reg}<22'b0101011011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011011000100000010) && ({row_reg, col_reg}<22'b0101011011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011011000100101101) && ({row_reg, col_reg}<22'b0101011011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011011001101010111) && ({row_reg, col_reg}<22'b0101011011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011011001110000010) && ({row_reg, col_reg}<22'b0101011011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011011010000000010) && ({row_reg, col_reg}<22'b0101011011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011011010000101101) && ({row_reg, col_reg}<22'b0101011011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011011100001010111) && ({row_reg, col_reg}<22'b0101011011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011011100010000010) && ({row_reg, col_reg}<22'b0101011011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011011100100000010) && ({row_reg, col_reg}<22'b0101011011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011011100100101101) && ({row_reg, col_reg}<22'b0101011011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011011101101010111) && ({row_reg, col_reg}<22'b0101011011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011011101110000010) && ({row_reg, col_reg}<22'b0101011011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011011110000000010) && ({row_reg, col_reg}<22'b0101011011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011011110000101101) && ({row_reg, col_reg}<22'b0101011100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011100000001010111) && ({row_reg, col_reg}<22'b0101011100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011100000010000010) && ({row_reg, col_reg}<22'b0101011100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011100000100000010) && ({row_reg, col_reg}<22'b0101011100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011100000100101101) && ({row_reg, col_reg}<22'b0101011100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011100001101010111) && ({row_reg, col_reg}<22'b0101011100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011100001110000010) && ({row_reg, col_reg}<22'b0101011100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011100010000000010) && ({row_reg, col_reg}<22'b0101011100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011100010000101101) && ({row_reg, col_reg}<22'b0101011100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011100100001010111) && ({row_reg, col_reg}<22'b0101011100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011100100010000010) && ({row_reg, col_reg}<22'b0101011100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011100100100000010) && ({row_reg, col_reg}<22'b0101011100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011100100100101101) && ({row_reg, col_reg}<22'b0101011100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011100101101010111) && ({row_reg, col_reg}<22'b0101011100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011100101110000010) && ({row_reg, col_reg}<22'b0101011100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011100110000000010) && ({row_reg, col_reg}<22'b0101011100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011100110000101101) && ({row_reg, col_reg}<22'b0101011101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011101000001010111) && ({row_reg, col_reg}<22'b0101011101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101011101000010000010) && ({row_reg, col_reg}<22'b0101011101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011101000100000010) && ({row_reg, col_reg}<22'b0101011101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011101000100101101) && ({row_reg, col_reg}<22'b0101011101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011101001101010111) && ({row_reg, col_reg}<22'b0101011101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011101001110000010) && ({row_reg, col_reg}<22'b0101011101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011101010000000010) && ({row_reg, col_reg}<22'b0101011101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011101010000101101) && ({row_reg, col_reg}<22'b0101011101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011101100001010111) && ({row_reg, col_reg}<22'b0101011101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101011101100010000010) && ({row_reg, col_reg}<22'b0101011101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011101100100000010) && ({row_reg, col_reg}<22'b0101011101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011101100100101101) && ({row_reg, col_reg}<22'b0101011101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011101101101010111) && ({row_reg, col_reg}<22'b0101011101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011101101110000010) && ({row_reg, col_reg}<22'b0101011101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011101110000000010) && ({row_reg, col_reg}<22'b0101011101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011101110000101101) && ({row_reg, col_reg}<22'b0101011110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011110000001010111) && ({row_reg, col_reg}<22'b0101011110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101011110000010000010) && ({row_reg, col_reg}<22'b0101011110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011110000100000010) && ({row_reg, col_reg}<22'b0101011110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011110000100101101) && ({row_reg, col_reg}<22'b0101011110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011110001101010111) && ({row_reg, col_reg}<22'b0101011110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011110001110000010) && ({row_reg, col_reg}<22'b0101011110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011110010000000010) && ({row_reg, col_reg}<22'b0101011110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011110010000101101) && ({row_reg, col_reg}<22'b0101011110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011110100001010111) && ({row_reg, col_reg}<22'b0101011110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011110100010000010) && ({row_reg, col_reg}<22'b0101011110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011110100100000010) && ({row_reg, col_reg}<22'b0101011110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011110100100101101) && ({row_reg, col_reg}<22'b0101011110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011110101101010111) && ({row_reg, col_reg}<22'b0101011110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011110101110000010) && ({row_reg, col_reg}<22'b0101011110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011110110000000010) && ({row_reg, col_reg}<22'b0101011110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011110110000101101) && ({row_reg, col_reg}<22'b0101011111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011111000001010111) && ({row_reg, col_reg}<22'b0101011111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101011111000010000010) && ({row_reg, col_reg}<22'b0101011111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011111000100000010) && ({row_reg, col_reg}<22'b0101011111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011111000100101101) && ({row_reg, col_reg}<22'b0101011111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011111001101010111) && ({row_reg, col_reg}<22'b0101011111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011111001110000010) && ({row_reg, col_reg}<22'b0101011111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011111010000000010) && ({row_reg, col_reg}<22'b0101011111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011111010000101101) && ({row_reg, col_reg}<22'b0101011111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011111100001010111) && ({row_reg, col_reg}<22'b0101011111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011111100010000010) && ({row_reg, col_reg}<22'b0101011111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011111100100000010) && ({row_reg, col_reg}<22'b0101011111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011111100100101101) && ({row_reg, col_reg}<22'b0101011111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101011111101101010111) && ({row_reg, col_reg}<22'b0101011111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101011111101110000010) && ({row_reg, col_reg}<22'b0101011111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101011111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101011111110000000010) && ({row_reg, col_reg}<22'b0101011111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101011111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101011111110000101101) && ({row_reg, col_reg}<22'b0101100000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100000000001010111) && ({row_reg, col_reg}<22'b0101100000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100000000010000010) && ({row_reg, col_reg}<22'b0101100000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100000000100000010) && ({row_reg, col_reg}<22'b0101100000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100000000100101101) && ({row_reg, col_reg}<22'b0101100000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100000001101010111) && ({row_reg, col_reg}<22'b0101100000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100000001110000010) && ({row_reg, col_reg}<22'b0101100000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100000010000000010) && ({row_reg, col_reg}<22'b0101100000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100000010000101101) && ({row_reg, col_reg}<22'b0101100000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100000100001010111) && ({row_reg, col_reg}<22'b0101100000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100000100010000010) && ({row_reg, col_reg}<22'b0101100000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100000100100000010) && ({row_reg, col_reg}<22'b0101100000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100000100100101101) && ({row_reg, col_reg}<22'b0101100000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100000101101010111) && ({row_reg, col_reg}<22'b0101100000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100000101110000010) && ({row_reg, col_reg}<22'b0101100000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100000110000000010) && ({row_reg, col_reg}<22'b0101100000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100000110000101101) && ({row_reg, col_reg}<22'b0101100001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100001000001010111) && ({row_reg, col_reg}<22'b0101100001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100001000010000010) && ({row_reg, col_reg}<22'b0101100001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100001000100000010) && ({row_reg, col_reg}<22'b0101100001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100001000100101101) && ({row_reg, col_reg}<22'b0101100001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100001001101010111) && ({row_reg, col_reg}<22'b0101100001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100001001110000010) && ({row_reg, col_reg}<22'b0101100001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100001010000000010) && ({row_reg, col_reg}<22'b0101100001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100001010000101101) && ({row_reg, col_reg}<22'b0101100001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100001100001010111) && ({row_reg, col_reg}<22'b0101100001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100001100010000010) && ({row_reg, col_reg}<22'b0101100001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100001100100000010) && ({row_reg, col_reg}<22'b0101100001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100001100100101101) && ({row_reg, col_reg}<22'b0101100001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100001101101010111) && ({row_reg, col_reg}<22'b0101100001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100001101110000010) && ({row_reg, col_reg}<22'b0101100001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100001110000000010) && ({row_reg, col_reg}<22'b0101100001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100001110000101101) && ({row_reg, col_reg}<22'b0101100010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100010000001010111) && ({row_reg, col_reg}<22'b0101100010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100010000010000010) && ({row_reg, col_reg}<22'b0101100010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100010000100000010) && ({row_reg, col_reg}<22'b0101100010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100010000100101101) && ({row_reg, col_reg}<22'b0101100010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100010001101010111) && ({row_reg, col_reg}<22'b0101100010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101100010001110000010) && ({row_reg, col_reg}<22'b0101100010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100010010000000010) && ({row_reg, col_reg}<22'b0101100010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100010010000101101) && ({row_reg, col_reg}<22'b0101100010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100010100001010111) && ({row_reg, col_reg}<22'b0101100010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100010100010000010) && ({row_reg, col_reg}<22'b0101100010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100010100100000010) && ({row_reg, col_reg}<22'b0101100010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100010100100101101) && ({row_reg, col_reg}<22'b0101100010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100010101101010111) && ({row_reg, col_reg}<22'b0101100010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101100010101110000010) && ({row_reg, col_reg}<22'b0101100010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100010110000000010) && ({row_reg, col_reg}<22'b0101100010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100010110000101101) && ({row_reg, col_reg}<22'b0101100011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100011000001010111) && ({row_reg, col_reg}<22'b0101100011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100011000010000010) && ({row_reg, col_reg}<22'b0101100011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100011000100000010) && ({row_reg, col_reg}<22'b0101100011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100011000100101101) && ({row_reg, col_reg}<22'b0101100011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100011001101010111) && ({row_reg, col_reg}<22'b0101100011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101100011001110000010) && ({row_reg, col_reg}<22'b0101100011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100011010000000010) && ({row_reg, col_reg}<22'b0101100011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100011010000101101) && ({row_reg, col_reg}<22'b0101100011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100011100001010111) && ({row_reg, col_reg}<22'b0101100011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100011100010000010) && ({row_reg, col_reg}<22'b0101100011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100011100100000010) && ({row_reg, col_reg}<22'b0101100011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100011100100101101) && ({row_reg, col_reg}<22'b0101100011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100011101101010111) && ({row_reg, col_reg}<22'b0101100011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101100011101110000010) && ({row_reg, col_reg}<22'b0101100011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100011110000000010) && ({row_reg, col_reg}<22'b0101100011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100011110000101101) && ({row_reg, col_reg}<22'b0101100100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100100000001010111) && ({row_reg, col_reg}<22'b0101100100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100100000010000010) && ({row_reg, col_reg}<22'b0101100100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100100000100000010) && ({row_reg, col_reg}<22'b0101100100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100100000100101101) && ({row_reg, col_reg}<22'b0101100100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100100001101010111) && ({row_reg, col_reg}<22'b0101100100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101100100001110000010) && ({row_reg, col_reg}<22'b0101100100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100100010000000010) && ({row_reg, col_reg}<22'b0101100100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100100010000101101) && ({row_reg, col_reg}<22'b0101100100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100100100001010111) && ({row_reg, col_reg}<22'b0101100100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100100100010000010) && ({row_reg, col_reg}<22'b0101100100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100100100100000010) && ({row_reg, col_reg}<22'b0101100100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100100100100101101) && ({row_reg, col_reg}<22'b0101100100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100100101101010111) && ({row_reg, col_reg}<22'b0101100100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101100100101110000010) && ({row_reg, col_reg}<22'b0101100100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100100110000000010) && ({row_reg, col_reg}<22'b0101100100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100100110000101101) && ({row_reg, col_reg}<22'b0101100101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100101000001010111) && ({row_reg, col_reg}<22'b0101100101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100101000010000010) && ({row_reg, col_reg}<22'b0101100101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100101000100000010) && ({row_reg, col_reg}<22'b0101100101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100101000100101101) && ({row_reg, col_reg}<22'b0101100101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100101001101010111) && ({row_reg, col_reg}<22'b0101100101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101100101001110000010) && ({row_reg, col_reg}<22'b0101100101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100101010000000010) && ({row_reg, col_reg}<22'b0101100101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100101010000101101) && ({row_reg, col_reg}<22'b0101100101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100101100001010111) && ({row_reg, col_reg}<22'b0101100101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100101100010000010) && ({row_reg, col_reg}<22'b0101100101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100101100100000010) && ({row_reg, col_reg}<22'b0101100101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100101100100101101) && ({row_reg, col_reg}<22'b0101100101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100101101101010111) && ({row_reg, col_reg}<22'b0101100101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100101101110000010) && ({row_reg, col_reg}<22'b0101100101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100101110000000010) && ({row_reg, col_reg}<22'b0101100101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100101110000101101) && ({row_reg, col_reg}<22'b0101100110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100110000001010111) && ({row_reg, col_reg}<22'b0101100110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101100110000010000010) && ({row_reg, col_reg}<22'b0101100110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100110000100000010) && ({row_reg, col_reg}<22'b0101100110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100110000100101101) && ({row_reg, col_reg}<22'b0101100110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100110001101010111) && ({row_reg, col_reg}<22'b0101100110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100110001110000010) && ({row_reg, col_reg}<22'b0101100110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100110010000000010) && ({row_reg, col_reg}<22'b0101100110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100110010000101101) && ({row_reg, col_reg}<22'b0101100110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100110100001010111) && ({row_reg, col_reg}<22'b0101100110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101100110100010000010) && ({row_reg, col_reg}<22'b0101100110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100110100100000010) && ({row_reg, col_reg}<22'b0101100110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100110100100101101) && ({row_reg, col_reg}<22'b0101100110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100110101101010111) && ({row_reg, col_reg}<22'b0101100110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100110101110000010) && ({row_reg, col_reg}<22'b0101100110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100110110000000010) && ({row_reg, col_reg}<22'b0101100110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100110110000101101) && ({row_reg, col_reg}<22'b0101100111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100111000001010111) && ({row_reg, col_reg}<22'b0101100111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101100111000010000010) && ({row_reg, col_reg}<22'b0101100111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100111000100000010) && ({row_reg, col_reg}<22'b0101100111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100111000100101101) && ({row_reg, col_reg}<22'b0101100111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100111001101010111) && ({row_reg, col_reg}<22'b0101100111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100111001110000010) && ({row_reg, col_reg}<22'b0101100111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100111010000000010) && ({row_reg, col_reg}<22'b0101100111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100111010000101101) && ({row_reg, col_reg}<22'b0101100111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100111100001010111) && ({row_reg, col_reg}<22'b0101100111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101100111100010000010) && ({row_reg, col_reg}<22'b0101100111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100111100100000010) && ({row_reg, col_reg}<22'b0101100111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100111100100101101) && ({row_reg, col_reg}<22'b0101100111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101100111101101010111) && ({row_reg, col_reg}<22'b0101100111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101100111101110000010) && ({row_reg, col_reg}<22'b0101100111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101100111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101100111110000000010) && ({row_reg, col_reg}<22'b0101100111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101100111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101100111110000101101) && ({row_reg, col_reg}<22'b0101101000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101000000001010111) && ({row_reg, col_reg}<22'b0101101000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101101000000010000010) && ({row_reg, col_reg}<22'b0101101000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101000000100000010) && ({row_reg, col_reg}<22'b0101101000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101000000100101101) && ({row_reg, col_reg}<22'b0101101000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101000001101010111) && ({row_reg, col_reg}<22'b0101101000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101000001110000010) && ({row_reg, col_reg}<22'b0101101000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101000010000000010) && ({row_reg, col_reg}<22'b0101101000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101000010000101101) && ({row_reg, col_reg}<22'b0101101000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101000100001010111) && ({row_reg, col_reg}<22'b0101101000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101101000100010000010) && ({row_reg, col_reg}<22'b0101101000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101000100100000010) && ({row_reg, col_reg}<22'b0101101000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101000100100101101) && ({row_reg, col_reg}<22'b0101101000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101000101101010111) && ({row_reg, col_reg}<22'b0101101000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101000101110000010) && ({row_reg, col_reg}<22'b0101101000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101000110000000010) && ({row_reg, col_reg}<22'b0101101000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101000110000101101) && ({row_reg, col_reg}<22'b0101101001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101001000001010111) && ({row_reg, col_reg}<22'b0101101001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101101001000010000010) && ({row_reg, col_reg}<22'b0101101001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101001000100000010) && ({row_reg, col_reg}<22'b0101101001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101001000100101101) && ({row_reg, col_reg}<22'b0101101001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101001001101010111) && ({row_reg, col_reg}<22'b0101101001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101001001110000010) && ({row_reg, col_reg}<22'b0101101001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101001010000000010) && ({row_reg, col_reg}<22'b0101101001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101001010000101101) && ({row_reg, col_reg}<22'b0101101001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101001100001010111) && ({row_reg, col_reg}<22'b0101101001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101001100010000010) && ({row_reg, col_reg}<22'b0101101001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101001100100000010) && ({row_reg, col_reg}<22'b0101101001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101001100100101101) && ({row_reg, col_reg}<22'b0101101001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101001101101010111) && ({row_reg, col_reg}<22'b0101101001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101001101110000010) && ({row_reg, col_reg}<22'b0101101001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101001110000000010) && ({row_reg, col_reg}<22'b0101101001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101001110000101101) && ({row_reg, col_reg}<22'b0101101010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101010000001010111) && ({row_reg, col_reg}<22'b0101101010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101010000010000010) && ({row_reg, col_reg}<22'b0101101010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101010000100000010) && ({row_reg, col_reg}<22'b0101101010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101010000100101101) && ({row_reg, col_reg}<22'b0101101010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101010001101010111) && ({row_reg, col_reg}<22'b0101101010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101010001110000010) && ({row_reg, col_reg}<22'b0101101010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101010010000000010) && ({row_reg, col_reg}<22'b0101101010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101010010000101101) && ({row_reg, col_reg}<22'b0101101010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101010100001010111) && ({row_reg, col_reg}<22'b0101101010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101010100010000010) && ({row_reg, col_reg}<22'b0101101010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101010100100000010) && ({row_reg, col_reg}<22'b0101101010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101010100100101101) && ({row_reg, col_reg}<22'b0101101010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101010101101010111) && ({row_reg, col_reg}<22'b0101101010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101010101110000010) && ({row_reg, col_reg}<22'b0101101010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101010110000000010) && ({row_reg, col_reg}<22'b0101101010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101010110000101101) && ({row_reg, col_reg}<22'b0101101011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101011000001010111) && ({row_reg, col_reg}<22'b0101101011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101011000010000010) && ({row_reg, col_reg}<22'b0101101011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101011000100000010) && ({row_reg, col_reg}<22'b0101101011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101011000100101101) && ({row_reg, col_reg}<22'b0101101011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101011001101010111) && ({row_reg, col_reg}<22'b0101101011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101011001110000010) && ({row_reg, col_reg}<22'b0101101011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101011010000000010) && ({row_reg, col_reg}<22'b0101101011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101011010000101101) && ({row_reg, col_reg}<22'b0101101011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101011100001010111) && ({row_reg, col_reg}<22'b0101101011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101011100010000010) && ({row_reg, col_reg}<22'b0101101011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101011100100000010) && ({row_reg, col_reg}<22'b0101101011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101011100100101101) && ({row_reg, col_reg}<22'b0101101011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101011101101010111) && ({row_reg, col_reg}<22'b0101101011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101011101110000010) && ({row_reg, col_reg}<22'b0101101011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101011110000000010) && ({row_reg, col_reg}<22'b0101101011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101011110000101101) && ({row_reg, col_reg}<22'b0101101100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101100000001010111) && ({row_reg, col_reg}<22'b0101101100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101100000010000010) && ({row_reg, col_reg}<22'b0101101100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101100000100000010) && ({row_reg, col_reg}<22'b0101101100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101100000100101101) && ({row_reg, col_reg}<22'b0101101100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101100001101010111) && ({row_reg, col_reg}<22'b0101101100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101101100001110000010) && ({row_reg, col_reg}<22'b0101101100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101100010000000010) && ({row_reg, col_reg}<22'b0101101100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101100010000101101) && ({row_reg, col_reg}<22'b0101101100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101100100001010111) && ({row_reg, col_reg}<22'b0101101100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101100100010000010) && ({row_reg, col_reg}<22'b0101101100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101100100100000010) && ({row_reg, col_reg}<22'b0101101100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101100100100101101) && ({row_reg, col_reg}<22'b0101101100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101100101101010111) && ({row_reg, col_reg}<22'b0101101100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101101100101110000010) && ({row_reg, col_reg}<22'b0101101100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101100110000000010) && ({row_reg, col_reg}<22'b0101101100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101100110000101101) && ({row_reg, col_reg}<22'b0101101101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101101000001010111) && ({row_reg, col_reg}<22'b0101101101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101101000010000010) && ({row_reg, col_reg}<22'b0101101101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101101000100000010) && ({row_reg, col_reg}<22'b0101101101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101101000100101101) && ({row_reg, col_reg}<22'b0101101101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101101001101010111) && ({row_reg, col_reg}<22'b0101101101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101101101001110000010) && ({row_reg, col_reg}<22'b0101101101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101101010000000010) && ({row_reg, col_reg}<22'b0101101101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101101010000101101) && ({row_reg, col_reg}<22'b0101101101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101101100001010111) && ({row_reg, col_reg}<22'b0101101101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101101100010000010) && ({row_reg, col_reg}<22'b0101101101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101101100100000010) && ({row_reg, col_reg}<22'b0101101101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101101100100101101) && ({row_reg, col_reg}<22'b0101101101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101101101101010111) && ({row_reg, col_reg}<22'b0101101101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101101101101110000010) && ({row_reg, col_reg}<22'b0101101101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101101110000000010) && ({row_reg, col_reg}<22'b0101101101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101101110000101101) && ({row_reg, col_reg}<22'b0101101110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101110000001010111) && ({row_reg, col_reg}<22'b0101101110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101110000010000010) && ({row_reg, col_reg}<22'b0101101110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101110000100000010) && ({row_reg, col_reg}<22'b0101101110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101110000100101101) && ({row_reg, col_reg}<22'b0101101110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101110001101010111) && ({row_reg, col_reg}<22'b0101101110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101101110001110000010) && ({row_reg, col_reg}<22'b0101101110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101110010000000010) && ({row_reg, col_reg}<22'b0101101110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101110010000101101) && ({row_reg, col_reg}<22'b0101101110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101110100001010111) && ({row_reg, col_reg}<22'b0101101110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101110100010000010) && ({row_reg, col_reg}<22'b0101101110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101110100100000010) && ({row_reg, col_reg}<22'b0101101110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101110100100101101) && ({row_reg, col_reg}<22'b0101101110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101110101101010111) && ({row_reg, col_reg}<22'b0101101110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101101110101110000010) && ({row_reg, col_reg}<22'b0101101110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101110110000000010) && ({row_reg, col_reg}<22'b0101101110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101110110000101101) && ({row_reg, col_reg}<22'b0101101111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101111000001010111) && ({row_reg, col_reg}<22'b0101101111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101111000010000010) && ({row_reg, col_reg}<22'b0101101111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101111000100000010) && ({row_reg, col_reg}<22'b0101101111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101111000100101101) && ({row_reg, col_reg}<22'b0101101111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101111001101010111) && ({row_reg, col_reg}<22'b0101101111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101101111001110000010) && ({row_reg, col_reg}<22'b0101101111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101111010000000010) && ({row_reg, col_reg}<22'b0101101111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101111010000101101) && ({row_reg, col_reg}<22'b0101101111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101111100001010111) && ({row_reg, col_reg}<22'b0101101111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101111100010000010) && ({row_reg, col_reg}<22'b0101101111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101111100100000010) && ({row_reg, col_reg}<22'b0101101111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101111100100101101) && ({row_reg, col_reg}<22'b0101101111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101101111101101010111) && ({row_reg, col_reg}<22'b0101101111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101101111101110000010) && ({row_reg, col_reg}<22'b0101101111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101101111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101101111110000000010) && ({row_reg, col_reg}<22'b0101101111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101101111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101101111110000101101) && ({row_reg, col_reg}<22'b0101110000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110000000001010111) && ({row_reg, col_reg}<22'b0101110000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101110000000010000010) && ({row_reg, col_reg}<22'b0101110000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110000000100000010) && ({row_reg, col_reg}<22'b0101110000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110000000100101101) && ({row_reg, col_reg}<22'b0101110000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110000001101010111) && ({row_reg, col_reg}<22'b0101110000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110000001110000010) && ({row_reg, col_reg}<22'b0101110000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110000010000000010) && ({row_reg, col_reg}<22'b0101110000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110000010000101101) && ({row_reg, col_reg}<22'b0101110000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110000100001010111) && ({row_reg, col_reg}<22'b0101110000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101110000100010000010) && ({row_reg, col_reg}<22'b0101110000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110000100100000010) && ({row_reg, col_reg}<22'b0101110000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110000100100101101) && ({row_reg, col_reg}<22'b0101110000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110000101101010111) && ({row_reg, col_reg}<22'b0101110000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110000101110000010) && ({row_reg, col_reg}<22'b0101110000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110000110000000010) && ({row_reg, col_reg}<22'b0101110000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110000110000101101) && ({row_reg, col_reg}<22'b0101110001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110001000001010111) && ({row_reg, col_reg}<22'b0101110001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101110001000010000010) && ({row_reg, col_reg}<22'b0101110001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110001000100000010) && ({row_reg, col_reg}<22'b0101110001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110001000100101101) && ({row_reg, col_reg}<22'b0101110001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110001001101010111) && ({row_reg, col_reg}<22'b0101110001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110001001110000010) && ({row_reg, col_reg}<22'b0101110001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110001010000000010) && ({row_reg, col_reg}<22'b0101110001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110001010000101101) && ({row_reg, col_reg}<22'b0101110001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110001100001010111) && ({row_reg, col_reg}<22'b0101110001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101110001100010000010) && ({row_reg, col_reg}<22'b0101110001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110001100100000010) && ({row_reg, col_reg}<22'b0101110001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110001100100101101) && ({row_reg, col_reg}<22'b0101110001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110001101101010111) && ({row_reg, col_reg}<22'b0101110001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110001101110000010) && ({row_reg, col_reg}<22'b0101110001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110001110000000010) && ({row_reg, col_reg}<22'b0101110001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110001110000101101) && ({row_reg, col_reg}<22'b0101110010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110010000001010111) && ({row_reg, col_reg}<22'b0101110010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101110010000010000010) && ({row_reg, col_reg}<22'b0101110010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110010000100000010) && ({row_reg, col_reg}<22'b0101110010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110010000100101101) && ({row_reg, col_reg}<22'b0101110010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110010001101010111) && ({row_reg, col_reg}<22'b0101110010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110010001110000010) && ({row_reg, col_reg}<22'b0101110010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110010010000000010) && ({row_reg, col_reg}<22'b0101110010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110010010000101101) && ({row_reg, col_reg}<22'b0101110010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110010100001010111) && ({row_reg, col_reg}<22'b0101110010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101110010100010000010) && ({row_reg, col_reg}<22'b0101110010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110010100100000010) && ({row_reg, col_reg}<22'b0101110010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110010100100101101) && ({row_reg, col_reg}<22'b0101110010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110010101101010111) && ({row_reg, col_reg}<22'b0101110010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110010101110000010) && ({row_reg, col_reg}<22'b0101110010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110010110000000010) && ({row_reg, col_reg}<22'b0101110010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110010110000101101) && ({row_reg, col_reg}<22'b0101110011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110011000001010111) && ({row_reg, col_reg}<22'b0101110011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101110011000010000010) && ({row_reg, col_reg}<22'b0101110011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110011000100000010) && ({row_reg, col_reg}<22'b0101110011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110011000100101101) && ({row_reg, col_reg}<22'b0101110011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110011001101010111) && ({row_reg, col_reg}<22'b0101110011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110011001110000010) && ({row_reg, col_reg}<22'b0101110011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110011010000000010) && ({row_reg, col_reg}<22'b0101110011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110011010000101101) && ({row_reg, col_reg}<22'b0101110011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110011100001010111) && ({row_reg, col_reg}<22'b0101110011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110011100010000010) && ({row_reg, col_reg}<22'b0101110011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110011100100000010) && ({row_reg, col_reg}<22'b0101110011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110011100100101101) && ({row_reg, col_reg}<22'b0101110011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110011101101010111) && ({row_reg, col_reg}<22'b0101110011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110011101110000010) && ({row_reg, col_reg}<22'b0101110011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110011110000000010) && ({row_reg, col_reg}<22'b0101110011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110011110000101101) && ({row_reg, col_reg}<22'b0101110100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110100000001010111) && ({row_reg, col_reg}<22'b0101110100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110100000010000010) && ({row_reg, col_reg}<22'b0101110100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110100000100000010) && ({row_reg, col_reg}<22'b0101110100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110100000100101101) && ({row_reg, col_reg}<22'b0101110100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110100001101010111) && ({row_reg, col_reg}<22'b0101110100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110100001110000010) && ({row_reg, col_reg}<22'b0101110100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110100010000000010) && ({row_reg, col_reg}<22'b0101110100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110100010000101101) && ({row_reg, col_reg}<22'b0101110100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110100100001010111) && ({row_reg, col_reg}<22'b0101110100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110100100010000010) && ({row_reg, col_reg}<22'b0101110100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110100100100000010) && ({row_reg, col_reg}<22'b0101110100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110100100100101101) && ({row_reg, col_reg}<22'b0101110100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110100101101010111) && ({row_reg, col_reg}<22'b0101110100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110100101110000010) && ({row_reg, col_reg}<22'b0101110100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110100110000000010) && ({row_reg, col_reg}<22'b0101110100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110100110000101101) && ({row_reg, col_reg}<22'b0101110101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110101000001010111) && ({row_reg, col_reg}<22'b0101110101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110101000010000010) && ({row_reg, col_reg}<22'b0101110101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110101000100000010) && ({row_reg, col_reg}<22'b0101110101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110101000100101101) && ({row_reg, col_reg}<22'b0101110101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110101001101010111) && ({row_reg, col_reg}<22'b0101110101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110101001110000010) && ({row_reg, col_reg}<22'b0101110101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110101010000000010) && ({row_reg, col_reg}<22'b0101110101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110101010000101101) && ({row_reg, col_reg}<22'b0101110101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110101100001010111) && ({row_reg, col_reg}<22'b0101110101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110101100010000010) && ({row_reg, col_reg}<22'b0101110101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110101100100000010) && ({row_reg, col_reg}<22'b0101110101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110101100100101101) && ({row_reg, col_reg}<22'b0101110101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110101101101010111) && ({row_reg, col_reg}<22'b0101110101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110101101110000010) && ({row_reg, col_reg}<22'b0101110101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110101110000000010) && ({row_reg, col_reg}<22'b0101110101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110101110000101101) && ({row_reg, col_reg}<22'b0101110110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110110000001010111) && ({row_reg, col_reg}<22'b0101110110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110110000010000010) && ({row_reg, col_reg}<22'b0101110110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110110000100000010) && ({row_reg, col_reg}<22'b0101110110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110110000100101101) && ({row_reg, col_reg}<22'b0101110110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110110001101010111) && ({row_reg, col_reg}<22'b0101110110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101110110001110000010) && ({row_reg, col_reg}<22'b0101110110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110110010000000010) && ({row_reg, col_reg}<22'b0101110110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110110010000101101) && ({row_reg, col_reg}<22'b0101110110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110110100001010111) && ({row_reg, col_reg}<22'b0101110110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110110100010000010) && ({row_reg, col_reg}<22'b0101110110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110110100100000010) && ({row_reg, col_reg}<22'b0101110110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110110100100101101) && ({row_reg, col_reg}<22'b0101110110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110110101101010111) && ({row_reg, col_reg}<22'b0101110110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101110110101110000010) && ({row_reg, col_reg}<22'b0101110110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110110110000000010) && ({row_reg, col_reg}<22'b0101110110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110110110000101101) && ({row_reg, col_reg}<22'b0101110111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110111000001010111) && ({row_reg, col_reg}<22'b0101110111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110111000010000010) && ({row_reg, col_reg}<22'b0101110111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110111000100000010) && ({row_reg, col_reg}<22'b0101110111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110111000100101101) && ({row_reg, col_reg}<22'b0101110111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110111001101010111) && ({row_reg, col_reg}<22'b0101110111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101110111001110000010) && ({row_reg, col_reg}<22'b0101110111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110111010000000010) && ({row_reg, col_reg}<22'b0101110111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110111010000101101) && ({row_reg, col_reg}<22'b0101110111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110111100001010111) && ({row_reg, col_reg}<22'b0101110111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101110111100010000010) && ({row_reg, col_reg}<22'b0101110111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110111100100000010) && ({row_reg, col_reg}<22'b0101110111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110111100100101101) && ({row_reg, col_reg}<22'b0101110111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101110111101101010111) && ({row_reg, col_reg}<22'b0101110111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101110111101110000010) && ({row_reg, col_reg}<22'b0101110111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101110111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101110111110000000010) && ({row_reg, col_reg}<22'b0101110111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101110111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101110111110000101101) && ({row_reg, col_reg}<22'b0101111000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111000000001010111) && ({row_reg, col_reg}<22'b0101111000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111000000010000010) && ({row_reg, col_reg}<22'b0101111000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111000000100000010) && ({row_reg, col_reg}<22'b0101111000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111000000100101101) && ({row_reg, col_reg}<22'b0101111000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111000001101010111) && ({row_reg, col_reg}<22'b0101111000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101111000001110000010) && ({row_reg, col_reg}<22'b0101111000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111000010000000010) && ({row_reg, col_reg}<22'b0101111000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111000010000101101) && ({row_reg, col_reg}<22'b0101111000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111000100001010111) && ({row_reg, col_reg}<22'b0101111000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111000100010000010) && ({row_reg, col_reg}<22'b0101111000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111000100100000010) && ({row_reg, col_reg}<22'b0101111000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111000100100101101) && ({row_reg, col_reg}<22'b0101111000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111000101101010111) && ({row_reg, col_reg}<22'b0101111000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101111000101110000010) && ({row_reg, col_reg}<22'b0101111000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111000110000000010) && ({row_reg, col_reg}<22'b0101111000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111000110000101101) && ({row_reg, col_reg}<22'b0101111001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111001000001010111) && ({row_reg, col_reg}<22'b0101111001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111001000010000010) && ({row_reg, col_reg}<22'b0101111001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111001000100000010) && ({row_reg, col_reg}<22'b0101111001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111001000100101101) && ({row_reg, col_reg}<22'b0101111001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111001001101010111) && ({row_reg, col_reg}<22'b0101111001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101111001001110000010) && ({row_reg, col_reg}<22'b0101111001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111001010000000010) && ({row_reg, col_reg}<22'b0101111001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111001010000101101) && ({row_reg, col_reg}<22'b0101111001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111001100001010111) && ({row_reg, col_reg}<22'b0101111001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111001100010000010) && ({row_reg, col_reg}<22'b0101111001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111001100100000010) && ({row_reg, col_reg}<22'b0101111001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111001100100101101) && ({row_reg, col_reg}<22'b0101111001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111001101101010111) && ({row_reg, col_reg}<22'b0101111001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111001101110000010) && ({row_reg, col_reg}<22'b0101111001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111001110000000010) && ({row_reg, col_reg}<22'b0101111001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111001110000101101) && ({row_reg, col_reg}<22'b0101111010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111010000001010111) && ({row_reg, col_reg}<22'b0101111010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101111010000010000010) && ({row_reg, col_reg}<22'b0101111010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111010000100000010) && ({row_reg, col_reg}<22'b0101111010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111010000100101101) && ({row_reg, col_reg}<22'b0101111010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111010001101010111) && ({row_reg, col_reg}<22'b0101111010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111010001110000010) && ({row_reg, col_reg}<22'b0101111010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111010010000000010) && ({row_reg, col_reg}<22'b0101111010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111010010000101101) && ({row_reg, col_reg}<22'b0101111010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111010100001010111) && ({row_reg, col_reg}<22'b0101111010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101111010100010000010) && ({row_reg, col_reg}<22'b0101111010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111010100100000010) && ({row_reg, col_reg}<22'b0101111010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111010100100101101) && ({row_reg, col_reg}<22'b0101111010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111010101101010111) && ({row_reg, col_reg}<22'b0101111010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111010101110000010) && ({row_reg, col_reg}<22'b0101111010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111010110000000010) && ({row_reg, col_reg}<22'b0101111010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111010110000101101) && ({row_reg, col_reg}<22'b0101111011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111011000001010111) && ({row_reg, col_reg}<22'b0101111011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101111011000010000010) && ({row_reg, col_reg}<22'b0101111011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111011000100000010) && ({row_reg, col_reg}<22'b0101111011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111011000100101101) && ({row_reg, col_reg}<22'b0101111011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111011001101010111) && ({row_reg, col_reg}<22'b0101111011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111011001110000010) && ({row_reg, col_reg}<22'b0101111011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111011010000000010) && ({row_reg, col_reg}<22'b0101111011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111011010000101101) && ({row_reg, col_reg}<22'b0101111011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111011100001010111) && ({row_reg, col_reg}<22'b0101111011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101111011100010000010) && ({row_reg, col_reg}<22'b0101111011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111011100100000010) && ({row_reg, col_reg}<22'b0101111011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111011100100101101) && ({row_reg, col_reg}<22'b0101111011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111011101101010111) && ({row_reg, col_reg}<22'b0101111011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111011101110000010) && ({row_reg, col_reg}<22'b0101111011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111011110000000010) && ({row_reg, col_reg}<22'b0101111011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111011110000101101) && ({row_reg, col_reg}<22'b0101111100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111100000001010111) && ({row_reg, col_reg}<22'b0101111100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0101111100000010000010) && ({row_reg, col_reg}<22'b0101111100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111100000100000010) && ({row_reg, col_reg}<22'b0101111100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111100000100101101) && ({row_reg, col_reg}<22'b0101111100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111100001101010111) && ({row_reg, col_reg}<22'b0101111100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111100001110000010) && ({row_reg, col_reg}<22'b0101111100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111100010000000010) && ({row_reg, col_reg}<22'b0101111100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111100010000101101) && ({row_reg, col_reg}<22'b0101111100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111100100001010111) && ({row_reg, col_reg}<22'b0101111100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101111100100010000010) && ({row_reg, col_reg}<22'b0101111100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111100100100000010) && ({row_reg, col_reg}<22'b0101111100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111100100100101101) && ({row_reg, col_reg}<22'b0101111100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111100101101010111) && ({row_reg, col_reg}<22'b0101111100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111100101110000010) && ({row_reg, col_reg}<22'b0101111100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111100110000000010) && ({row_reg, col_reg}<22'b0101111100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111100110000101101) && ({row_reg, col_reg}<22'b0101111101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111101000001010111) && ({row_reg, col_reg}<22'b0101111101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0101111101000010000010) && ({row_reg, col_reg}<22'b0101111101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111101000100000010) && ({row_reg, col_reg}<22'b0101111101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111101000100101101) && ({row_reg, col_reg}<22'b0101111101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111101001101010111) && ({row_reg, col_reg}<22'b0101111101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111101001110000010) && ({row_reg, col_reg}<22'b0101111101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111101010000000010) && ({row_reg, col_reg}<22'b0101111101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111101010000101101) && ({row_reg, col_reg}<22'b0101111101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111101100001010111) && ({row_reg, col_reg}<22'b0101111101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111101100010000010) && ({row_reg, col_reg}<22'b0101111101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111101100100000010) && ({row_reg, col_reg}<22'b0101111101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111101100100101101) && ({row_reg, col_reg}<22'b0101111101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111101101101010111) && ({row_reg, col_reg}<22'b0101111101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111101101110000010) && ({row_reg, col_reg}<22'b0101111101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111101110000000010) && ({row_reg, col_reg}<22'b0101111101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111101110000101101) && ({row_reg, col_reg}<22'b0101111110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111110000001010111) && ({row_reg, col_reg}<22'b0101111110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111110000010000010) && ({row_reg, col_reg}<22'b0101111110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111110000100000010) && ({row_reg, col_reg}<22'b0101111110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111110000100101101) && ({row_reg, col_reg}<22'b0101111110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111110001101010111) && ({row_reg, col_reg}<22'b0101111110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111110001110000010) && ({row_reg, col_reg}<22'b0101111110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111110010000000010) && ({row_reg, col_reg}<22'b0101111110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111110010000101101) && ({row_reg, col_reg}<22'b0101111110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111110100001010111) && ({row_reg, col_reg}<22'b0101111110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111110100010000010) && ({row_reg, col_reg}<22'b0101111110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111110100100000010) && ({row_reg, col_reg}<22'b0101111110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111110100100101101) && ({row_reg, col_reg}<22'b0101111110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111110101101010111) && ({row_reg, col_reg}<22'b0101111110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111110101110000010) && ({row_reg, col_reg}<22'b0101111110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111110110000000010) && ({row_reg, col_reg}<22'b0101111110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111110110000101101) && ({row_reg, col_reg}<22'b0101111111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111111000001010111) && ({row_reg, col_reg}<22'b0101111111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111111000010000010) && ({row_reg, col_reg}<22'b0101111111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111111000100000010) && ({row_reg, col_reg}<22'b0101111111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111111000100101101) && ({row_reg, col_reg}<22'b0101111111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111111001101010111) && ({row_reg, col_reg}<22'b0101111111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111111001110000010) && ({row_reg, col_reg}<22'b0101111111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111111010000000010) && ({row_reg, col_reg}<22'b0101111111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111111010000101101) && ({row_reg, col_reg}<22'b0101111111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111111100001010111) && ({row_reg, col_reg}<22'b0101111111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111111100010000010) && ({row_reg, col_reg}<22'b0101111111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111111100100000010) && ({row_reg, col_reg}<22'b0101111111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111111100100101101) && ({row_reg, col_reg}<22'b0101111111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0101111111101101010111) && ({row_reg, col_reg}<22'b0101111111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0101111111101110000010) && ({row_reg, col_reg}<22'b0101111111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0101111111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0101111111110000000010) && ({row_reg, col_reg}<22'b0101111111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0101111111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0101111111110000101101) && ({row_reg, col_reg}<22'b0110000000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000000000001010111) && ({row_reg, col_reg}<22'b0110000000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000000000010000010) && ({row_reg, col_reg}<22'b0110000000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000000000100000010) && ({row_reg, col_reg}<22'b0110000000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000000000100101101) && ({row_reg, col_reg}<22'b0110000000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000000001101010111) && ({row_reg, col_reg}<22'b0110000000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000000001110000010) && ({row_reg, col_reg}<22'b0110000000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000000010000000010) && ({row_reg, col_reg}<22'b0110000000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000000010000101101) && ({row_reg, col_reg}<22'b0110000000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000000100001010111) && ({row_reg, col_reg}<22'b0110000000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000000100010000010) && ({row_reg, col_reg}<22'b0110000000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000000100100000010) && ({row_reg, col_reg}<22'b0110000000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000000100100101101) && ({row_reg, col_reg}<22'b0110000000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000000101101010111) && ({row_reg, col_reg}<22'b0110000000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000000101110000010) && ({row_reg, col_reg}<22'b0110000000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000000110000000010) && ({row_reg, col_reg}<22'b0110000000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000000110000101101) && ({row_reg, col_reg}<22'b0110000001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000001000001010111) && ({row_reg, col_reg}<22'b0110000001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000001000010000010) && ({row_reg, col_reg}<22'b0110000001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000001000100000010) && ({row_reg, col_reg}<22'b0110000001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000001000100101101) && ({row_reg, col_reg}<22'b0110000001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000001001101010111) && ({row_reg, col_reg}<22'b0110000001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110000001001110000010) && ({row_reg, col_reg}<22'b0110000001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000001010000000010) && ({row_reg, col_reg}<22'b0110000001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000001010000101101) && ({row_reg, col_reg}<22'b0110000001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000001100001010111) && ({row_reg, col_reg}<22'b0110000001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000001100010000010) && ({row_reg, col_reg}<22'b0110000001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000001100100000010) && ({row_reg, col_reg}<22'b0110000001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000001100100101101) && ({row_reg, col_reg}<22'b0110000001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000001101101010111) && ({row_reg, col_reg}<22'b0110000001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110000001101110000010) && ({row_reg, col_reg}<22'b0110000001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000001110000000010) && ({row_reg, col_reg}<22'b0110000001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000001110000101101) && ({row_reg, col_reg}<22'b0110000010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000010000001010111) && ({row_reg, col_reg}<22'b0110000010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000010000010000010) && ({row_reg, col_reg}<22'b0110000010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000010000100000010) && ({row_reg, col_reg}<22'b0110000010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000010000100101101) && ({row_reg, col_reg}<22'b0110000010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000010001101010111) && ({row_reg, col_reg}<22'b0110000010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110000010001110000010) && ({row_reg, col_reg}<22'b0110000010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000010010000000010) && ({row_reg, col_reg}<22'b0110000010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000010010000101101) && ({row_reg, col_reg}<22'b0110000010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000010100001010111) && ({row_reg, col_reg}<22'b0110000010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000010100010000010) && ({row_reg, col_reg}<22'b0110000010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000010100100000010) && ({row_reg, col_reg}<22'b0110000010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000010100100101101) && ({row_reg, col_reg}<22'b0110000010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000010101101010111) && ({row_reg, col_reg}<22'b0110000010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000010101110000010) && ({row_reg, col_reg}<22'b0110000010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000010110000000010) && ({row_reg, col_reg}<22'b0110000010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000010110000101101) && ({row_reg, col_reg}<22'b0110000011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000011000001010111) && ({row_reg, col_reg}<22'b0110000011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000011000010000010) && ({row_reg, col_reg}<22'b0110000011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000011000100000010) && ({row_reg, col_reg}<22'b0110000011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000011000100101101) && ({row_reg, col_reg}<22'b0110000011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000011001101010111) && ({row_reg, col_reg}<22'b0110000011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000011001110000010) && ({row_reg, col_reg}<22'b0110000011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000011010000000010) && ({row_reg, col_reg}<22'b0110000011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000011010000101101) && ({row_reg, col_reg}<22'b0110000011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000011100001010111) && ({row_reg, col_reg}<22'b0110000011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000011100010000010) && ({row_reg, col_reg}<22'b0110000011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000011100100000010) && ({row_reg, col_reg}<22'b0110000011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000011100100101101) && ({row_reg, col_reg}<22'b0110000011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000011101101010111) && ({row_reg, col_reg}<22'b0110000011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000011101110000010) && ({row_reg, col_reg}<22'b0110000011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000011110000000010) && ({row_reg, col_reg}<22'b0110000011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000011110000101101) && ({row_reg, col_reg}<22'b0110000100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000100000001010111) && ({row_reg, col_reg}<22'b0110000100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000100000010000010) && ({row_reg, col_reg}<22'b0110000100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000100000100000010) && ({row_reg, col_reg}<22'b0110000100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000100000100101101) && ({row_reg, col_reg}<22'b0110000100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000100001101010111) && ({row_reg, col_reg}<22'b0110000100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000100001110000010) && ({row_reg, col_reg}<22'b0110000100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000100010000000010) && ({row_reg, col_reg}<22'b0110000100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000100010000101101) && ({row_reg, col_reg}<22'b0110000100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000100100001010111) && ({row_reg, col_reg}<22'b0110000100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000100100010000010) && ({row_reg, col_reg}<22'b0110000100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000100100100000010) && ({row_reg, col_reg}<22'b0110000100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000100100100101101) && ({row_reg, col_reg}<22'b0110000100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000100101101010111) && ({row_reg, col_reg}<22'b0110000100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000100101110000010) && ({row_reg, col_reg}<22'b0110000100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000100110000000010) && ({row_reg, col_reg}<22'b0110000100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000100110000101101) && ({row_reg, col_reg}<22'b0110000101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000101000001010111) && ({row_reg, col_reg}<22'b0110000101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110000101000010000010) && ({row_reg, col_reg}<22'b0110000101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000101000100000010) && ({row_reg, col_reg}<22'b0110000101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000101000100101101) && ({row_reg, col_reg}<22'b0110000101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000101001101010111) && ({row_reg, col_reg}<22'b0110000101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000101001110000010) && ({row_reg, col_reg}<22'b0110000101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000101010000000010) && ({row_reg, col_reg}<22'b0110000101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000101010000101101) && ({row_reg, col_reg}<22'b0110000101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000101100001010111) && ({row_reg, col_reg}<22'b0110000101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110000101100010000010) && ({row_reg, col_reg}<22'b0110000101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000101100100000010) && ({row_reg, col_reg}<22'b0110000101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000101100100101101) && ({row_reg, col_reg}<22'b0110000101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000101101101010111) && ({row_reg, col_reg}<22'b0110000101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000101101110000010) && ({row_reg, col_reg}<22'b0110000101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000101110000000010) && ({row_reg, col_reg}<22'b0110000101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000101110000101101) && ({row_reg, col_reg}<22'b0110000110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000110000001010111) && ({row_reg, col_reg}<22'b0110000110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110000110000010000010) && ({row_reg, col_reg}<22'b0110000110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000110000100000010) && ({row_reg, col_reg}<22'b0110000110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000110000100101101) && ({row_reg, col_reg}<22'b0110000110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000110001101010111) && ({row_reg, col_reg}<22'b0110000110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000110001110000010) && ({row_reg, col_reg}<22'b0110000110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000110010000000010) && ({row_reg, col_reg}<22'b0110000110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000110010000101101) && ({row_reg, col_reg}<22'b0110000110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000110100001010111) && ({row_reg, col_reg}<22'b0110000110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000110100010000010) && ({row_reg, col_reg}<22'b0110000110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000110100100000010) && ({row_reg, col_reg}<22'b0110000110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000110100100101101) && ({row_reg, col_reg}<22'b0110000110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000110101101010111) && ({row_reg, col_reg}<22'b0110000110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000110101110000010) && ({row_reg, col_reg}<22'b0110000110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000110110000000010) && ({row_reg, col_reg}<22'b0110000110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000110110000101101) && ({row_reg, col_reg}<22'b0110000111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000111000001010111) && ({row_reg, col_reg}<22'b0110000111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110000111000010000010) && ({row_reg, col_reg}<22'b0110000111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000111000100000010) && ({row_reg, col_reg}<22'b0110000111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000111000100101101) && ({row_reg, col_reg}<22'b0110000111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000111001101010111) && ({row_reg, col_reg}<22'b0110000111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000111001110000010) && ({row_reg, col_reg}<22'b0110000111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000111010000000010) && ({row_reg, col_reg}<22'b0110000111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000111010000101101) && ({row_reg, col_reg}<22'b0110000111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000111100001010111) && ({row_reg, col_reg}<22'b0110000111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000111100010000010) && ({row_reg, col_reg}<22'b0110000111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000111100100000010) && ({row_reg, col_reg}<22'b0110000111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000111100100101101) && ({row_reg, col_reg}<22'b0110000111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110000111101101010111) && ({row_reg, col_reg}<22'b0110000111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110000111101110000010) && ({row_reg, col_reg}<22'b0110000111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110000111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110000111110000000010) && ({row_reg, col_reg}<22'b0110000111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110000111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110000111110000101101) && ({row_reg, col_reg}<22'b0110001000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001000000001010111) && ({row_reg, col_reg}<22'b0110001000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001000000010000010) && ({row_reg, col_reg}<22'b0110001000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001000000100000010) && ({row_reg, col_reg}<22'b0110001000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001000000100101101) && ({row_reg, col_reg}<22'b0110001000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001000001101010111) && ({row_reg, col_reg}<22'b0110001000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001000001110000010) && ({row_reg, col_reg}<22'b0110001000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001000010000000010) && ({row_reg, col_reg}<22'b0110001000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001000010000101101) && ({row_reg, col_reg}<22'b0110001000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001000100001010111) && ({row_reg, col_reg}<22'b0110001000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001000100010000010) && ({row_reg, col_reg}<22'b0110001000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001000100100000010) && ({row_reg, col_reg}<22'b0110001000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001000100100101101) && ({row_reg, col_reg}<22'b0110001000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001000101101010111) && ({row_reg, col_reg}<22'b0110001000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001000101110000010) && ({row_reg, col_reg}<22'b0110001000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001000110000000010) && ({row_reg, col_reg}<22'b0110001000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001000110000101101) && ({row_reg, col_reg}<22'b0110001001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001001000001010111) && ({row_reg, col_reg}<22'b0110001001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001001000010000010) && ({row_reg, col_reg}<22'b0110001001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001001000100000010) && ({row_reg, col_reg}<22'b0110001001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001001000100101101) && ({row_reg, col_reg}<22'b0110001001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001001001101010111) && ({row_reg, col_reg}<22'b0110001001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001001001110000010) && ({row_reg, col_reg}<22'b0110001001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001001010000000010) && ({row_reg, col_reg}<22'b0110001001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001001010000101101) && ({row_reg, col_reg}<22'b0110001001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001001100001010111) && ({row_reg, col_reg}<22'b0110001001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001001100010000010) && ({row_reg, col_reg}<22'b0110001001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001001100100000010) && ({row_reg, col_reg}<22'b0110001001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001001100100101101) && ({row_reg, col_reg}<22'b0110001001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001001101101010111) && ({row_reg, col_reg}<22'b0110001001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001001101110000010) && ({row_reg, col_reg}<22'b0110001001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001001110000000010) && ({row_reg, col_reg}<22'b0110001001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001001110000101101) && ({row_reg, col_reg}<22'b0110001010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001010000001010111) && ({row_reg, col_reg}<22'b0110001010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001010000010000010) && ({row_reg, col_reg}<22'b0110001010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001010000100000010) && ({row_reg, col_reg}<22'b0110001010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001010000100101101) && ({row_reg, col_reg}<22'b0110001010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001010001101010111) && ({row_reg, col_reg}<22'b0110001010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110001010001110000010) && ({row_reg, col_reg}<22'b0110001010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001010010000000010) && ({row_reg, col_reg}<22'b0110001010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001010010000101101) && ({row_reg, col_reg}<22'b0110001010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001010100001010111) && ({row_reg, col_reg}<22'b0110001010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001010100010000010) && ({row_reg, col_reg}<22'b0110001010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001010100100000010) && ({row_reg, col_reg}<22'b0110001010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001010100100101101) && ({row_reg, col_reg}<22'b0110001010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001010101101010111) && ({row_reg, col_reg}<22'b0110001010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110001010101110000010) && ({row_reg, col_reg}<22'b0110001010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001010110000000010) && ({row_reg, col_reg}<22'b0110001010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001010110000101101) && ({row_reg, col_reg}<22'b0110001011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001011000001010111) && ({row_reg, col_reg}<22'b0110001011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001011000010000010) && ({row_reg, col_reg}<22'b0110001011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001011000100000010) && ({row_reg, col_reg}<22'b0110001011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001011000100101101) && ({row_reg, col_reg}<22'b0110001011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001011001101010111) && ({row_reg, col_reg}<22'b0110001011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110001011001110000010) && ({row_reg, col_reg}<22'b0110001011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001011010000000010) && ({row_reg, col_reg}<22'b0110001011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001011010000101101) && ({row_reg, col_reg}<22'b0110001011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001011100001010111) && ({row_reg, col_reg}<22'b0110001011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001011100010000010) && ({row_reg, col_reg}<22'b0110001011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001011100100000010) && ({row_reg, col_reg}<22'b0110001011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001011100100101101) && ({row_reg, col_reg}<22'b0110001011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001011101101010111) && ({row_reg, col_reg}<22'b0110001011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110001011101110000010) && ({row_reg, col_reg}<22'b0110001011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001011110000000010) && ({row_reg, col_reg}<22'b0110001011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001011110000101101) && ({row_reg, col_reg}<22'b0110001100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001100000001010111) && ({row_reg, col_reg}<22'b0110001100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001100000010000010) && ({row_reg, col_reg}<22'b0110001100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001100000100000010) && ({row_reg, col_reg}<22'b0110001100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001100000100101101) && ({row_reg, col_reg}<22'b0110001100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001100001101010111) && ({row_reg, col_reg}<22'b0110001100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110001100001110000010) && ({row_reg, col_reg}<22'b0110001100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001100010000000010) && ({row_reg, col_reg}<22'b0110001100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001100010000101101) && ({row_reg, col_reg}<22'b0110001100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001100100001010111) && ({row_reg, col_reg}<22'b0110001100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001100100010000010) && ({row_reg, col_reg}<22'b0110001100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001100100100000010) && ({row_reg, col_reg}<22'b0110001100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001100100100101101) && ({row_reg, col_reg}<22'b0110001100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001100101101010111) && ({row_reg, col_reg}<22'b0110001100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110001100101110000010) && ({row_reg, col_reg}<22'b0110001100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001100110000000010) && ({row_reg, col_reg}<22'b0110001100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001100110000101101) && ({row_reg, col_reg}<22'b0110001101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001101000001010111) && ({row_reg, col_reg}<22'b0110001101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001101000010000010) && ({row_reg, col_reg}<22'b0110001101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001101000100000010) && ({row_reg, col_reg}<22'b0110001101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001101000100101101) && ({row_reg, col_reg}<22'b0110001101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001101001101010111) && ({row_reg, col_reg}<22'b0110001101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110001101001110000010) && ({row_reg, col_reg}<22'b0110001101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001101010000000010) && ({row_reg, col_reg}<22'b0110001101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001101010000101101) && ({row_reg, col_reg}<22'b0110001101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001101100001010111) && ({row_reg, col_reg}<22'b0110001101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001101100010000010) && ({row_reg, col_reg}<22'b0110001101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001101100100000010) && ({row_reg, col_reg}<22'b0110001101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001101100100101101) && ({row_reg, col_reg}<22'b0110001101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001101101101010111) && ({row_reg, col_reg}<22'b0110001101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001101101110000010) && ({row_reg, col_reg}<22'b0110001101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001101110000000010) && ({row_reg, col_reg}<22'b0110001101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001101110000101101) && ({row_reg, col_reg}<22'b0110001110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001110000001010111) && ({row_reg, col_reg}<22'b0110001110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110001110000010000010) && ({row_reg, col_reg}<22'b0110001110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001110000100000010) && ({row_reg, col_reg}<22'b0110001110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001110000100101101) && ({row_reg, col_reg}<22'b0110001110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001110001101010111) && ({row_reg, col_reg}<22'b0110001110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001110001110000010) && ({row_reg, col_reg}<22'b0110001110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001110010000000010) && ({row_reg, col_reg}<22'b0110001110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001110010000101101) && ({row_reg, col_reg}<22'b0110001110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001110100001010111) && ({row_reg, col_reg}<22'b0110001110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110001110100010000010) && ({row_reg, col_reg}<22'b0110001110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001110100100000010) && ({row_reg, col_reg}<22'b0110001110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001110100100101101) && ({row_reg, col_reg}<22'b0110001110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001110101101010111) && ({row_reg, col_reg}<22'b0110001110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001110101110000010) && ({row_reg, col_reg}<22'b0110001110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001110110000000010) && ({row_reg, col_reg}<22'b0110001110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001110110000101101) && ({row_reg, col_reg}<22'b0110001111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001111000001010111) && ({row_reg, col_reg}<22'b0110001111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110001111000010000010) && ({row_reg, col_reg}<22'b0110001111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001111000100000010) && ({row_reg, col_reg}<22'b0110001111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001111000100101101) && ({row_reg, col_reg}<22'b0110001111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001111001101010111) && ({row_reg, col_reg}<22'b0110001111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001111001110000010) && ({row_reg, col_reg}<22'b0110001111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001111010000000010) && ({row_reg, col_reg}<22'b0110001111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001111010000101101) && ({row_reg, col_reg}<22'b0110001111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001111100001010111) && ({row_reg, col_reg}<22'b0110001111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110001111100010000010) && ({row_reg, col_reg}<22'b0110001111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001111100100000010) && ({row_reg, col_reg}<22'b0110001111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001111100100101101) && ({row_reg, col_reg}<22'b0110001111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110001111101101010111) && ({row_reg, col_reg}<22'b0110001111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110001111101110000010) && ({row_reg, col_reg}<22'b0110001111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110001111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110001111110000000010) && ({row_reg, col_reg}<22'b0110001111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110001111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110001111110000101101) && ({row_reg, col_reg}<22'b0110010000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010000000001010111) && ({row_reg, col_reg}<22'b0110010000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110010000000010000010) && ({row_reg, col_reg}<22'b0110010000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010000000100000010) && ({row_reg, col_reg}<22'b0110010000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010000000100101101) && ({row_reg, col_reg}<22'b0110010000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010000001101010111) && ({row_reg, col_reg}<22'b0110010000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010000001110000010) && ({row_reg, col_reg}<22'b0110010000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010000010000000010) && ({row_reg, col_reg}<22'b0110010000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010000010000101101) && ({row_reg, col_reg}<22'b0110010000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010000100001010111) && ({row_reg, col_reg}<22'b0110010000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110010000100010000010) && ({row_reg, col_reg}<22'b0110010000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010000100100000010) && ({row_reg, col_reg}<22'b0110010000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010000100100101101) && ({row_reg, col_reg}<22'b0110010000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010000101101010111) && ({row_reg, col_reg}<22'b0110010000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010000101110000010) && ({row_reg, col_reg}<22'b0110010000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010000110000000010) && ({row_reg, col_reg}<22'b0110010000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010000110000101101) && ({row_reg, col_reg}<22'b0110010001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010001000001010111) && ({row_reg, col_reg}<22'b0110010001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110010001000010000010) && ({row_reg, col_reg}<22'b0110010001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010001000100000010) && ({row_reg, col_reg}<22'b0110010001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010001000100101101) && ({row_reg, col_reg}<22'b0110010001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010001001101010111) && ({row_reg, col_reg}<22'b0110010001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010001001110000010) && ({row_reg, col_reg}<22'b0110010001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010001010000000010) && ({row_reg, col_reg}<22'b0110010001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010001010000101101) && ({row_reg, col_reg}<22'b0110010001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010001100001010111) && ({row_reg, col_reg}<22'b0110010001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010001100010000010) && ({row_reg, col_reg}<22'b0110010001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010001100100000010) && ({row_reg, col_reg}<22'b0110010001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010001100100101101) && ({row_reg, col_reg}<22'b0110010001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010001101101010111) && ({row_reg, col_reg}<22'b0110010001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010001101110000010) && ({row_reg, col_reg}<22'b0110010001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010001110000000010) && ({row_reg, col_reg}<22'b0110010001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010001110000101101) && ({row_reg, col_reg}<22'b0110010010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010010000001010111) && ({row_reg, col_reg}<22'b0110010010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010010000010000010) && ({row_reg, col_reg}<22'b0110010010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010010000100000010) && ({row_reg, col_reg}<22'b0110010010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010010000100101101) && ({row_reg, col_reg}<22'b0110010010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010010001101010111) && ({row_reg, col_reg}<22'b0110010010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010010001110000010) && ({row_reg, col_reg}<22'b0110010010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010010010000000010) && ({row_reg, col_reg}<22'b0110010010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010010010000101101) && ({row_reg, col_reg}<22'b0110010010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010010100001010111) && ({row_reg, col_reg}<22'b0110010010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010010100010000010) && ({row_reg, col_reg}<22'b0110010010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010010100100000010) && ({row_reg, col_reg}<22'b0110010010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010010100100101101) && ({row_reg, col_reg}<22'b0110010010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010010101101010111) && ({row_reg, col_reg}<22'b0110010010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010010101110000010) && ({row_reg, col_reg}<22'b0110010010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010010110000000010) && ({row_reg, col_reg}<22'b0110010010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010010110000101101) && ({row_reg, col_reg}<22'b0110010011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010011000001010111) && ({row_reg, col_reg}<22'b0110010011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010011000010000010) && ({row_reg, col_reg}<22'b0110010011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010011000100000010) && ({row_reg, col_reg}<22'b0110010011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010011000100101101) && ({row_reg, col_reg}<22'b0110010011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010011001101010111) && ({row_reg, col_reg}<22'b0110010011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010011001110000010) && ({row_reg, col_reg}<22'b0110010011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010011010000000010) && ({row_reg, col_reg}<22'b0110010011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010011010000101101) && ({row_reg, col_reg}<22'b0110010011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010011100001010111) && ({row_reg, col_reg}<22'b0110010011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010011100010000010) && ({row_reg, col_reg}<22'b0110010011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010011100100000010) && ({row_reg, col_reg}<22'b0110010011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010011100100101101) && ({row_reg, col_reg}<22'b0110010011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010011101101010111) && ({row_reg, col_reg}<22'b0110010011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010011101110000010) && ({row_reg, col_reg}<22'b0110010011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010011110000000010) && ({row_reg, col_reg}<22'b0110010011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010011110000101101) && ({row_reg, col_reg}<22'b0110010100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010100000001010111) && ({row_reg, col_reg}<22'b0110010100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010100000010000010) && ({row_reg, col_reg}<22'b0110010100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010100000100000010) && ({row_reg, col_reg}<22'b0110010100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010100000100101101) && ({row_reg, col_reg}<22'b0110010100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010100001101010111) && ({row_reg, col_reg}<22'b0110010100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110010100001110000010) && ({row_reg, col_reg}<22'b0110010100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010100010000000010) && ({row_reg, col_reg}<22'b0110010100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010100010000101101) && ({row_reg, col_reg}<22'b0110010100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010100100001010111) && ({row_reg, col_reg}<22'b0110010100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010100100010000010) && ({row_reg, col_reg}<22'b0110010100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010100100100000010) && ({row_reg, col_reg}<22'b0110010100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010100100100101101) && ({row_reg, col_reg}<22'b0110010100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010100101101010111) && ({row_reg, col_reg}<22'b0110010100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110010100101110000010) && ({row_reg, col_reg}<22'b0110010100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010100110000000010) && ({row_reg, col_reg}<22'b0110010100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010100110000101101) && ({row_reg, col_reg}<22'b0110010101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010101000001010111) && ({row_reg, col_reg}<22'b0110010101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010101000010000010) && ({row_reg, col_reg}<22'b0110010101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010101000100000010) && ({row_reg, col_reg}<22'b0110010101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010101000100101101) && ({row_reg, col_reg}<22'b0110010101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010101001101010111) && ({row_reg, col_reg}<22'b0110010101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110010101001110000010) && ({row_reg, col_reg}<22'b0110010101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010101010000000010) && ({row_reg, col_reg}<22'b0110010101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010101010000101101) && ({row_reg, col_reg}<22'b0110010101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010101100001010111) && ({row_reg, col_reg}<22'b0110010101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010101100010000010) && ({row_reg, col_reg}<22'b0110010101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010101100100000010) && ({row_reg, col_reg}<22'b0110010101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010101100100101101) && ({row_reg, col_reg}<22'b0110010101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010101101101010111) && ({row_reg, col_reg}<22'b0110010101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110010101101110000010) && ({row_reg, col_reg}<22'b0110010101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010101110000000010) && ({row_reg, col_reg}<22'b0110010101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010101110000101101) && ({row_reg, col_reg}<22'b0110010110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010110000001010111) && ({row_reg, col_reg}<22'b0110010110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010110000010000010) && ({row_reg, col_reg}<22'b0110010110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010110000100000010) && ({row_reg, col_reg}<22'b0110010110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010110000100101101) && ({row_reg, col_reg}<22'b0110010110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010110001101010111) && ({row_reg, col_reg}<22'b0110010110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110010110001110000010) && ({row_reg, col_reg}<22'b0110010110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010110010000000010) && ({row_reg, col_reg}<22'b0110010110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010110010000101101) && ({row_reg, col_reg}<22'b0110010110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010110100001010111) && ({row_reg, col_reg}<22'b0110010110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010110100010000010) && ({row_reg, col_reg}<22'b0110010110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010110100100000010) && ({row_reg, col_reg}<22'b0110010110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010110100100101101) && ({row_reg, col_reg}<22'b0110010110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010110101101010111) && ({row_reg, col_reg}<22'b0110010110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110010110101110000010) && ({row_reg, col_reg}<22'b0110010110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010110110000000010) && ({row_reg, col_reg}<22'b0110010110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010110110000101101) && ({row_reg, col_reg}<22'b0110010111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010111000001010111) && ({row_reg, col_reg}<22'b0110010111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010111000010000010) && ({row_reg, col_reg}<22'b0110010111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010111000100000010) && ({row_reg, col_reg}<22'b0110010111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010111000100101101) && ({row_reg, col_reg}<22'b0110010111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010111001101010111) && ({row_reg, col_reg}<22'b0110010111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110010111001110000010) && ({row_reg, col_reg}<22'b0110010111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010111010000000010) && ({row_reg, col_reg}<22'b0110010111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010111010000101101) && ({row_reg, col_reg}<22'b0110010111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010111100001010111) && ({row_reg, col_reg}<22'b0110010111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010111100010000010) && ({row_reg, col_reg}<22'b0110010111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010111100100000010) && ({row_reg, col_reg}<22'b0110010111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010111100100101101) && ({row_reg, col_reg}<22'b0110010111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110010111101101010111) && ({row_reg, col_reg}<22'b0110010111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110010111101110000010) && ({row_reg, col_reg}<22'b0110010111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110010111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110010111110000000010) && ({row_reg, col_reg}<22'b0110010111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110010111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110010111110000101101) && ({row_reg, col_reg}<22'b0110011000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011000000001010111) && ({row_reg, col_reg}<22'b0110011000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110011000000010000010) && ({row_reg, col_reg}<22'b0110011000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011000000100000010) && ({row_reg, col_reg}<22'b0110011000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011000000100101101) && ({row_reg, col_reg}<22'b0110011000001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011000001101010111) && ({row_reg, col_reg}<22'b0110011000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011000001110000010) && ({row_reg, col_reg}<22'b0110011000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011000010000000010) && ({row_reg, col_reg}<22'b0110011000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011000010000101101) && ({row_reg, col_reg}<22'b0110011000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011000100001010111) && ({row_reg, col_reg}<22'b0110011000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110011000100010000010) && ({row_reg, col_reg}<22'b0110011000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011000100100000010) && ({row_reg, col_reg}<22'b0110011000100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011000100100101101) && ({row_reg, col_reg}<22'b0110011000101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011000101101010111) && ({row_reg, col_reg}<22'b0110011000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011000101110000010) && ({row_reg, col_reg}<22'b0110011000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011000110000000010) && ({row_reg, col_reg}<22'b0110011000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011000110000101101) && ({row_reg, col_reg}<22'b0110011001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011001000001010111) && ({row_reg, col_reg}<22'b0110011001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110011001000010000010) && ({row_reg, col_reg}<22'b0110011001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011001000100000010) && ({row_reg, col_reg}<22'b0110011001000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011001000100101101) && ({row_reg, col_reg}<22'b0110011001001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011001001101010111) && ({row_reg, col_reg}<22'b0110011001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011001001110000010) && ({row_reg, col_reg}<22'b0110011001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011001010000000010) && ({row_reg, col_reg}<22'b0110011001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011001010000101101) && ({row_reg, col_reg}<22'b0110011001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011001100001010111) && ({row_reg, col_reg}<22'b0110011001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110011001100010000010) && ({row_reg, col_reg}<22'b0110011001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011001100100000010) && ({row_reg, col_reg}<22'b0110011001100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011001100100101101) && ({row_reg, col_reg}<22'b0110011001101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011001101101010111) && ({row_reg, col_reg}<22'b0110011001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011001101110000010) && ({row_reg, col_reg}<22'b0110011001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011001110000000010) && ({row_reg, col_reg}<22'b0110011001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011001110000101101) && ({row_reg, col_reg}<22'b0110011010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011010000001010111) && ({row_reg, col_reg}<22'b0110011010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110011010000010000010) && ({row_reg, col_reg}<22'b0110011010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011010000100000010) && ({row_reg, col_reg}<22'b0110011010000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011010000100101101) && ({row_reg, col_reg}<22'b0110011010001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011010001101010111) && ({row_reg, col_reg}<22'b0110011010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011010001110000010) && ({row_reg, col_reg}<22'b0110011010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011010010000000010) && ({row_reg, col_reg}<22'b0110011010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011010010000101101) && ({row_reg, col_reg}<22'b0110011010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011010100001010111) && ({row_reg, col_reg}<22'b0110011010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110011010100010000010) && ({row_reg, col_reg}<22'b0110011010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011010100100000010) && ({row_reg, col_reg}<22'b0110011010100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011010100100101101) && ({row_reg, col_reg}<22'b0110011010101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011010101101010111) && ({row_reg, col_reg}<22'b0110011010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011010101110000010) && ({row_reg, col_reg}<22'b0110011010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011010110000000010) && ({row_reg, col_reg}<22'b0110011010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011010110000101101) && ({row_reg, col_reg}<22'b0110011011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011011000001010111) && ({row_reg, col_reg}<22'b0110011011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110011011000010000010) && ({row_reg, col_reg}<22'b0110011011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011011000100000010) && ({row_reg, col_reg}<22'b0110011011000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011011000100101101) && ({row_reg, col_reg}<22'b0110011011001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011011001101010111) && ({row_reg, col_reg}<22'b0110011011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011011001110000010) && ({row_reg, col_reg}<22'b0110011011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011011010000000010) && ({row_reg, col_reg}<22'b0110011011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011011010000101101) && ({row_reg, col_reg}<22'b0110011011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011011100001010111) && ({row_reg, col_reg}<22'b0110011011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011011100010000010) && ({row_reg, col_reg}<22'b0110011011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011011100100000010) && ({row_reg, col_reg}<22'b0110011011100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011011100100101101) && ({row_reg, col_reg}<22'b0110011011101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011011101101010111) && ({row_reg, col_reg}<22'b0110011011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011011101110000010) && ({row_reg, col_reg}<22'b0110011011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011011110000000010) && ({row_reg, col_reg}<22'b0110011011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011011110000101101) && ({row_reg, col_reg}<22'b0110011100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011100000001010111) && ({row_reg, col_reg}<22'b0110011100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011100000010000010) && ({row_reg, col_reg}<22'b0110011100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011100000100000010) && ({row_reg, col_reg}<22'b0110011100000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011100000100101101) && ({row_reg, col_reg}<22'b0110011100001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011100001101010111) && ({row_reg, col_reg}<22'b0110011100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011100001110000010) && ({row_reg, col_reg}<22'b0110011100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011100010000000010) && ({row_reg, col_reg}<22'b0110011100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011100010000101101) && ({row_reg, col_reg}<22'b0110011100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011100100001010111) && ({row_reg, col_reg}<22'b0110011100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011100100010000010) && ({row_reg, col_reg}<22'b0110011100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011100100100000010) && ({row_reg, col_reg}<22'b0110011100100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011100100100101101) && ({row_reg, col_reg}<22'b0110011100101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011100101101010111) && ({row_reg, col_reg}<22'b0110011100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011100101110000010) && ({row_reg, col_reg}<22'b0110011100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011100110000000010) && ({row_reg, col_reg}<22'b0110011100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011100110000101101) && ({row_reg, col_reg}<22'b0110011101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011101000001010111) && ({row_reg, col_reg}<22'b0110011101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011101000010000010) && ({row_reg, col_reg}<22'b0110011101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011101000100000010) && ({row_reg, col_reg}<22'b0110011101000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011101000100101101) && ({row_reg, col_reg}<22'b0110011101001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011101001101010111) && ({row_reg, col_reg}<22'b0110011101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011101001110000010) && ({row_reg, col_reg}<22'b0110011101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011101010000000010) && ({row_reg, col_reg}<22'b0110011101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011101010000101101) && ({row_reg, col_reg}<22'b0110011101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011101100001010111) && ({row_reg, col_reg}<22'b0110011101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011101100010000010) && ({row_reg, col_reg}<22'b0110011101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011101100100000010) && ({row_reg, col_reg}<22'b0110011101100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011101100100101101) && ({row_reg, col_reg}<22'b0110011101101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011101101101010111) && ({row_reg, col_reg}<22'b0110011101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011101101110000010) && ({row_reg, col_reg}<22'b0110011101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011101110000000010) && ({row_reg, col_reg}<22'b0110011101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011101110000101101) && ({row_reg, col_reg}<22'b0110011110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011110000001010111) && ({row_reg, col_reg}<22'b0110011110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011110000010000010) && ({row_reg, col_reg}<22'b0110011110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011110000100000010) && ({row_reg, col_reg}<22'b0110011110000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011110000100101101) && ({row_reg, col_reg}<22'b0110011110001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011110001101010111) && ({row_reg, col_reg}<22'b0110011110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110011110001110000010) && ({row_reg, col_reg}<22'b0110011110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011110010000000010) && ({row_reg, col_reg}<22'b0110011110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011110010000101101) && ({row_reg, col_reg}<22'b0110011110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011110100001010111) && ({row_reg, col_reg}<22'b0110011110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011110100010000010) && ({row_reg, col_reg}<22'b0110011110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011110100100000010) && ({row_reg, col_reg}<22'b0110011110100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011110100100101101) && ({row_reg, col_reg}<22'b0110011110101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011110101101010111) && ({row_reg, col_reg}<22'b0110011110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110011110101110000010) && ({row_reg, col_reg}<22'b0110011110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011110110000000010) && ({row_reg, col_reg}<22'b0110011110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011110110000101101) && ({row_reg, col_reg}<22'b0110011111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011111000001010111) && ({row_reg, col_reg}<22'b0110011111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011111000010000010) && ({row_reg, col_reg}<22'b0110011111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011111000100000010) && ({row_reg, col_reg}<22'b0110011111000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111000100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011111000100101101) && ({row_reg, col_reg}<22'b0110011111001101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011111001101010111) && ({row_reg, col_reg}<22'b0110011111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110011111001110000010) && ({row_reg, col_reg}<22'b0110011111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011111010000000010) && ({row_reg, col_reg}<22'b0110011111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011111010000101101) && ({row_reg, col_reg}<22'b0110011111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011111100001010111) && ({row_reg, col_reg}<22'b0110011111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110011111100010000010) && ({row_reg, col_reg}<22'b0110011111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011111100100000010) && ({row_reg, col_reg}<22'b0110011111100100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111100100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011111100100101101) && ({row_reg, col_reg}<22'b0110011111101101010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110011111101101010111) && ({row_reg, col_reg}<22'b0110011111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110011111101110000010) && ({row_reg, col_reg}<22'b0110011111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110011111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110011111110000000010) && ({row_reg, col_reg}<22'b0110011111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110011111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110011111110000101101) && ({row_reg, col_reg}<22'b0110100000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100000000001010111) && ({row_reg, col_reg}<22'b0110100000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100000000010000010) && ({row_reg, col_reg}<22'b0110100000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100000000100000010) && ({row_reg, col_reg}<22'b0110100000000100101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000000100101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100000000100101101) && ({row_reg, col_reg}<22'b0110100000000111101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100000000111101101) && ({row_reg, col_reg}<22'b0110100000001010010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100000001010010110) && ({row_reg, col_reg}<22'b0110100000001101010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100000001101010111) && ({row_reg, col_reg}<22'b0110100000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110100000001110000010) && ({row_reg, col_reg}<22'b0110100000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100000010000000010) && ({row_reg, col_reg}<22'b0110100000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100000010000101101) && ({row_reg, col_reg}<22'b0110100000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100000100001010111) && ({row_reg, col_reg}<22'b0110100000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100000100010000010) && ({row_reg, col_reg}<22'b0110100000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100000100100000010) && ({row_reg, col_reg}<22'b0110100000100111110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000100111110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b0110100000100111110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0110100000100111110011) && ({row_reg, col_reg}<22'b0110100000101010010000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100000101010010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==22'b0110100000101010010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b0110100000101010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110100000101010010011) && ({row_reg, col_reg}<22'b0110100000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110100000101110000010) && ({row_reg, col_reg}<22'b0110100000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100000110000000010) && ({row_reg, col_reg}<22'b0110100000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100000110000101101) && ({row_reg, col_reg}<22'b0110100001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100001000001010111) && ({row_reg, col_reg}<22'b0110100001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100001000010000010) && ({row_reg, col_reg}<22'b0110100001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100001000100000010) && ({row_reg, col_reg}<22'b0110100001000111110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001000111110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0110100001000111110101) && ({row_reg, col_reg}<22'b0110100001001010001110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100001001010001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100001001010001111) && ({row_reg, col_reg}<22'b0110100001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110100001001110000010) && ({row_reg, col_reg}<22'b0110100001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100001010000000010) && ({row_reg, col_reg}<22'b0110100001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100001010000101101) && ({row_reg, col_reg}<22'b0110100001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100001100001010111) && ({row_reg, col_reg}<22'b0110100001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100001100010000010) && ({row_reg, col_reg}<22'b0110100001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100001100100000010) && ({row_reg, col_reg}<22'b0110100001100111110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001100111110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0110100001100111110111) && ({row_reg, col_reg}<22'b0110100001101010001100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100001101010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100001101010001101) && ({row_reg, col_reg}<22'b0110100001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100001101110000010) && ({row_reg, col_reg}<22'b0110100001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100001110000000010) && ({row_reg, col_reg}<22'b0110100001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100001110000101101) && ({row_reg, col_reg}<22'b0110100010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100010000001010111) && ({row_reg, col_reg}<22'b0110100010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110100010000010000010) && ({row_reg, col_reg}<22'b0110100010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100010000100000010) && ({row_reg, col_reg}<22'b0110100010000111111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010000111111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100010000111111001) && ({row_reg, col_reg}<22'b0110100010001010001011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100010001010001011) && ({row_reg, col_reg}<22'b0110100010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100010001110000010) && ({row_reg, col_reg}<22'b0110100010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100010010000000010) && ({row_reg, col_reg}<22'b0110100010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100010010000101101) && ({row_reg, col_reg}<22'b0110100010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100010100001010111) && ({row_reg, col_reg}<22'b0110100010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110100010100010000010) && ({row_reg, col_reg}<22'b0110100010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100010100100000010) && ({row_reg, col_reg}<22'b0110100010100111111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010100111111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0110100010100111111010) && ({row_reg, col_reg}<22'b0110100010101010001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100010101010001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100010101010001010) && ({row_reg, col_reg}<22'b0110100010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100010101110000010) && ({row_reg, col_reg}<22'b0110100010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100010110000000010) && ({row_reg, col_reg}<22'b0110100010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100010110000101101) && ({row_reg, col_reg}<22'b0110100011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100011000001010111) && ({row_reg, col_reg}<22'b0110100011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110100011000010000010) && ({row_reg, col_reg}<22'b0110100011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100011000100000010) && ({row_reg, col_reg}<22'b0110100011000111111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011000111111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110100011000111111011) && ({row_reg, col_reg}<22'b0110100011001010001000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100011001010001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100011001010001001) && ({row_reg, col_reg}<22'b0110100011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100011001110000010) && ({row_reg, col_reg}<22'b0110100011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100011010000000010) && ({row_reg, col_reg}<22'b0110100011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100011010000101101) && ({row_reg, col_reg}<22'b0110100011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100011100001010111) && ({row_reg, col_reg}<22'b0110100011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110100011100010000010) && ({row_reg, col_reg}<22'b0110100011100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100011100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100011100100000010) && ({row_reg, col_reg}<22'b0110100011100111111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011100111111011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0110100011100111111100) && ({row_reg, col_reg}<22'b0110100011101010000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100011101010000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100011101010001000) && ({row_reg, col_reg}<22'b0110100011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100011101110000010) && ({row_reg, col_reg}<22'b0110100011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100011110000000010) && ({row_reg, col_reg}<22'b0110100011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100011110000101101) && ({row_reg, col_reg}<22'b0110100100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100100000001010111) && ({row_reg, col_reg}<22'b0110100100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110100100000010000010) && ({row_reg, col_reg}<22'b0110100100000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100100000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100100000100000010) && ({row_reg, col_reg}<22'b0110100100000111111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100000111111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110100100000111111101) && ({row_reg, col_reg}<22'b0110100100001010000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100100001010000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100100001010000111) && ({row_reg, col_reg}<22'b0110100100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100100001110000010) && ({row_reg, col_reg}<22'b0110100100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100100010000000010) && ({row_reg, col_reg}<22'b0110100100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100100010000101101) && ({row_reg, col_reg}<22'b0110100100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100100100001010111) && ({row_reg, col_reg}<22'b0110100100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110100100100010000010) && ({row_reg, col_reg}<22'b0110100100100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100100100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100100100100000010) && ({row_reg, col_reg}<22'b0110100100100111111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100100111111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100100100111111110) && ({row_reg, col_reg}<22'b0110100100101010000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100100101010000110) && ({row_reg, col_reg}<22'b0110100100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100100101110000010) && ({row_reg, col_reg}<22'b0110100100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100100110000000010) && ({row_reg, col_reg}<22'b0110100100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100100110000101101) && ({row_reg, col_reg}<22'b0110100101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100101000001010111) && ({row_reg, col_reg}<22'b0110100101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110100101000010000010) && ({row_reg, col_reg}<22'b0110100101000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100101000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100101000100000010) && ({row_reg, col_reg}<22'b0110100101000111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110100101000111111110) && ({row_reg, col_reg}<22'b0110100101001010000101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100101001010000101) && ({row_reg, col_reg}<22'b0110100101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100101001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100101001110000010) && ({row_reg, col_reg}<22'b0110100101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100101010000000010) && ({row_reg, col_reg}<22'b0110100101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100101010000101101) && ({row_reg, col_reg}<22'b0110100101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100101100001010111) && ({row_reg, col_reg}<22'b0110100101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100101100010000010) && ({row_reg, col_reg}<22'b0110100101100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100101100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100101100100000010) && ({row_reg, col_reg}<22'b0110100101100111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100101100111111110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=22'b0110100101100111111111) && ({row_reg, col_reg}<22'b0110100101101010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100101101010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100101101010000101) && ({row_reg, col_reg}<22'b0110100101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100101101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100101101110000010) && ({row_reg, col_reg}<22'b0110100101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100101110000000010) && ({row_reg, col_reg}<22'b0110100101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100101110000101101) && ({row_reg, col_reg}<22'b0110100110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100110000001010111) && ({row_reg, col_reg}<22'b0110100110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100110000010000010) && ({row_reg, col_reg}<22'b0110100110000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100110000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100110000100000010) && ({row_reg, col_reg}<22'b0110100110000111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110000111111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0110100110001000000000) && ({row_reg, col_reg}<22'b0110100110001010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100110001010000100) && ({row_reg, col_reg}<22'b0110100110001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100110001110000010) && ({row_reg, col_reg}<22'b0110100110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100110010000000010) && ({row_reg, col_reg}<22'b0110100110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100110010000101101) && ({row_reg, col_reg}<22'b0110100110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100110100001010111) && ({row_reg, col_reg}<22'b0110100110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100110100010000010) && ({row_reg, col_reg}<22'b0110100110100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100110100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100110100100000010) && ({row_reg, col_reg}<22'b0110100110100111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110100111111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0110100110101000000000) && ({row_reg, col_reg}<22'b0110100110101010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100110101010000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110100110101010000100) && ({row_reg, col_reg}<22'b0110100110101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100110101110000010) && ({row_reg, col_reg}<22'b0110100110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100110110000000010) && ({row_reg, col_reg}<22'b0110100110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100110110000101101) && ({row_reg, col_reg}<22'b0110100111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100111000001010111) && ({row_reg, col_reg}<22'b0110100111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100111000010000010) && ({row_reg, col_reg}<22'b0110100111000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100111000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100111000100000010) && ({row_reg, col_reg}<22'b0110100111001000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110100111001000000000) && ({row_reg, col_reg}<22'b0110100111001010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100111001010000011) && ({row_reg, col_reg}<22'b0110100111001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100111001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100111001110000010) && ({row_reg, col_reg}<22'b0110100111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100111010000000010) && ({row_reg, col_reg}<22'b0110100111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100111010000101101) && ({row_reg, col_reg}<22'b0110100111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110100111100001010111) && ({row_reg, col_reg}<22'b0110100111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100111100010000010) && ({row_reg, col_reg}<22'b0110100111100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100111100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100111100100000010) && ({row_reg, col_reg}<22'b0110100111101000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100111101000000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100111101000000001) && ({row_reg, col_reg}<22'b0110100111101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100111101010000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100111101010000011) && ({row_reg, col_reg}<22'b0110100111101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100111101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110100111101110000010) && ({row_reg, col_reg}<22'b0110100111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110100111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110100111110000000010) && ({row_reg, col_reg}<22'b0110100111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110100111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110100111110000101101) && ({row_reg, col_reg}<22'b0110101000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101000000001010111) && ({row_reg, col_reg}<22'b0110101000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101000000010000010) && ({row_reg, col_reg}<22'b0110101000000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101000000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101000000100000010) && ({row_reg, col_reg}<22'b0110101000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110101000001000000001) && ({row_reg, col_reg}<22'b0110101000001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101000001010000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101000001010000011) && ({row_reg, col_reg}<22'b0110101000001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101000001110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101000001110000010) && ({row_reg, col_reg}<22'b0110101000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101000010000000010) && ({row_reg, col_reg}<22'b0110101000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101000010000101101) && ({row_reg, col_reg}<22'b0110101000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101000100001010111) && ({row_reg, col_reg}<22'b0110101000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101000100010000010) && ({row_reg, col_reg}<22'b0110101000100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101000100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101000100100000010) && ({row_reg, col_reg}<22'b0110101000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110101000101000000001) && ({row_reg, col_reg}<22'b0110101000101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101000101010000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110101000101010000011) && ({row_reg, col_reg}<22'b0110101000101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101000101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101000101110000010) && ({row_reg, col_reg}<22'b0110101000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101000110000000010) && ({row_reg, col_reg}<22'b0110101000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101000110000101101) && ({row_reg, col_reg}<22'b0110101001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101001000001010111) && ({row_reg, col_reg}<22'b0110101001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101001000010000010) && ({row_reg, col_reg}<22'b0110101001000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101001000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101001000100000010) && ({row_reg, col_reg}<22'b0110101001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001001000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101001001000000010) && ({row_reg, col_reg}<22'b0110101001001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101001001010000010) && ({row_reg, col_reg}<22'b0110101001001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101001001110000010) && ({row_reg, col_reg}<22'b0110101001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101001010000000010) && ({row_reg, col_reg}<22'b0110101001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101001010000101101) && ({row_reg, col_reg}<22'b0110101001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101001100001010111) && ({row_reg, col_reg}<22'b0110101001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101001100010000010) && ({row_reg, col_reg}<22'b0110101001100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101001100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101001100100000010) && ({row_reg, col_reg}<22'b0110101001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001101000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110101001101000000010) && ({row_reg, col_reg}<22'b0110101001101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101001101010000010) && ({row_reg, col_reg}<22'b0110101001101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001101110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101001101110000010) && ({row_reg, col_reg}<22'b0110101001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101001110000000010) && ({row_reg, col_reg}<22'b0110101001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101001110000101101) && ({row_reg, col_reg}<22'b0110101010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101010000001010111) && ({row_reg, col_reg}<22'b0110101010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101010000010000010) && ({row_reg, col_reg}<22'b0110101010000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101010000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101010000100000010) && ({row_reg, col_reg}<22'b0110101010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101010001000000010) && ({row_reg, col_reg}<22'b0110101010001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101010001010000010) && ({row_reg, col_reg}<22'b0110101010001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010001110000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101010001110000010) && ({row_reg, col_reg}<22'b0110101010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101010010000000010) && ({row_reg, col_reg}<22'b0110101010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101010010000101101) && ({row_reg, col_reg}<22'b0110101010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101010100001010111) && ({row_reg, col_reg}<22'b0110101010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101010100010000010) && ({row_reg, col_reg}<22'b0110101010100100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101010100100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101010100100000010) && ({row_reg, col_reg}<22'b0110101010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101010101000000010) && ({row_reg, col_reg}<22'b0110101010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101010101010000010) && ({row_reg, col_reg}<22'b0110101010101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010101110000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101010101110000010) && ({row_reg, col_reg}<22'b0110101010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101010110000000010) && ({row_reg, col_reg}<22'b0110101010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101010110000101101) && ({row_reg, col_reg}<22'b0110101011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101011000001010111) && ({row_reg, col_reg}<22'b0110101011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101011000010000010) && ({row_reg, col_reg}<22'b0110101011000100000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101011000100000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101011000100000010) && ({row_reg, col_reg}<22'b0110101011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101011001000000010) && ({row_reg, col_reg}<22'b0110101011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101011001010000010) && ({row_reg, col_reg}<22'b0110101011001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011001110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101011001110000010) && ({row_reg, col_reg}<22'b0110101011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101011010000000010) && ({row_reg, col_reg}<22'b0110101011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101011010000101101) && ({row_reg, col_reg}<22'b0110101011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101011100001010111) && ({row_reg, col_reg}<22'b0110101011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101011100010000010) && ({row_reg, col_reg}<22'b0110101011100100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101011100100000010) && ({row_reg, col_reg}<22'b0110101011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101011101000000010) && ({row_reg, col_reg}<22'b0110101011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101011101010000010) && ({row_reg, col_reg}<22'b0110101011101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011101110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101011101110000010) && ({row_reg, col_reg}<22'b0110101011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101011110000000010) && ({row_reg, col_reg}<22'b0110101011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101011110000101101) && ({row_reg, col_reg}<22'b0110101100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101100000001010111) && ({row_reg, col_reg}<22'b0110101100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101100000010000010) && ({row_reg, col_reg}<22'b0110101100000100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101100000100000010) && ({row_reg, col_reg}<22'b0110101100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101100001000000010) && ({row_reg, col_reg}<22'b0110101100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101100001010000010) && ({row_reg, col_reg}<22'b0110101100001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100001110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110101100001110000010) && ({row_reg, col_reg}<22'b0110101100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101100010000000010) && ({row_reg, col_reg}<22'b0110101100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101100010000101101) && ({row_reg, col_reg}<22'b0110101100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101100100001010111) && ({row_reg, col_reg}<22'b0110101100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101100100010000010) && ({row_reg, col_reg}<22'b0110101100100100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101100100100000010) && ({row_reg, col_reg}<22'b0110101100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101100101000000010) && ({row_reg, col_reg}<22'b0110101100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101100101010000010) && ({row_reg, col_reg}<22'b0110101100101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100101110000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101100101110000010) && ({row_reg, col_reg}<22'b0110101100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101100110000000010) && ({row_reg, col_reg}<22'b0110101100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101100110000101101) && ({row_reg, col_reg}<22'b0110101101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101101000001010111) && ({row_reg, col_reg}<22'b0110101101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101101000010000010) && ({row_reg, col_reg}<22'b0110101101000100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101101000100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110101101000100000011) && ({row_reg, col_reg}<22'b0110101101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101101001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101101001000000010) && ({row_reg, col_reg}<22'b0110101101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101101001010000010) && ({row_reg, col_reg}<22'b0110101101001110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110101101001110000001) && ({row_reg, col_reg}<22'b0110101101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101101010000000010) && ({row_reg, col_reg}<22'b0110101101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101101010000101101) && ({row_reg, col_reg}<22'b0110101101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101101100001010111) && ({row_reg, col_reg}<22'b0110101101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101101100010000010) && ({row_reg, col_reg}<22'b0110101101100100000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101101100100000011) && ({row_reg, col_reg}<22'b0110101101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101101101000000010) && ({row_reg, col_reg}<22'b0110101101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101101101010000010) && ({row_reg, col_reg}<22'b0110101101101110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110101101101110000001) && ({row_reg, col_reg}<22'b0110101101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101101110000000010) && ({row_reg, col_reg}<22'b0110101101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101101110000101101) && ({row_reg, col_reg}<22'b0110101110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101110000001010111) && ({row_reg, col_reg}<22'b0110101110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110101110000010000010) && ({row_reg, col_reg}<22'b0110101110000100000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101110000100000011) && ({row_reg, col_reg}<22'b0110101110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101110001000000010) && ({row_reg, col_reg}<22'b0110101110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101110001010000010) && ({row_reg, col_reg}<22'b0110101110001110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101110001110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101110001110000001) && ({row_reg, col_reg}<22'b0110101110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101110010000000010) && ({row_reg, col_reg}<22'b0110101110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101110010000101101) && ({row_reg, col_reg}<22'b0110101110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101110100001010111) && ({row_reg, col_reg}<22'b0110101110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101110100010000010) && ({row_reg, col_reg}<22'b0110101110100100000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101110100100000011) && ({row_reg, col_reg}<22'b0110101110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101110101000000010) && ({row_reg, col_reg}<22'b0110101110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101110101010000010) && ({row_reg, col_reg}<22'b0110101110101110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110101110101110000000) && ({row_reg, col_reg}<22'b0110101110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101110110000000010) && ({row_reg, col_reg}<22'b0110101110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101110110000101101) && ({row_reg, col_reg}<22'b0110101111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101111000001010111) && ({row_reg, col_reg}<22'b0110101111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110101111000010000010) && ({row_reg, col_reg}<22'b0110101111000100000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101111000100000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110101111000100000100) && ({row_reg, col_reg}<22'b0110101111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101111001000000010) && ({row_reg, col_reg}<22'b0110101111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101111001010000010) && ({row_reg, col_reg}<22'b0110101111001101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111001101111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0110101111001110000000) && ({row_reg, col_reg}<22'b0110101111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101111010000000010) && ({row_reg, col_reg}<22'b0110101111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101111010000101101) && ({row_reg, col_reg}<22'b0110101111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101111100001010111) && ({row_reg, col_reg}<22'b0110101111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101111100010000010) && ({row_reg, col_reg}<22'b0110101111100100000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110101111100100000100) && ({row_reg, col_reg}<22'b0110101111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110101111101000000010) && ({row_reg, col_reg}<22'b0110101111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101111101010000010) && ({row_reg, col_reg}<22'b0110101111101101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111101101111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0110101111101110000000) && ({row_reg, col_reg}<22'b0110101111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110101111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110101111110000000010) && ({row_reg, col_reg}<22'b0110101111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110101111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110101111110000101101) && ({row_reg, col_reg}<22'b0110110000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110000000001010111) && ({row_reg, col_reg}<22'b0110110000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110000000010000010) && ({row_reg, col_reg}<22'b0110110000000100000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110000000100000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110110000000100000101) && ({row_reg, col_reg}<22'b0110110000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110000001000000010) && ({row_reg, col_reg}<22'b0110110000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110000001010000010) && ({row_reg, col_reg}<22'b0110110000001101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110000001101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110110000001101111111) && ({row_reg, col_reg}<22'b0110110000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110000010000000010) && ({row_reg, col_reg}<22'b0110110000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110000010000101101) && ({row_reg, col_reg}<22'b0110110000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110000100001010111) && ({row_reg, col_reg}<22'b0110110000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110000100010000010) && ({row_reg, col_reg}<22'b0110110000100100000101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110000100100000101) && ({row_reg, col_reg}<22'b0110110000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110000101000000010) && ({row_reg, col_reg}<22'b0110110000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110000101010000010) && ({row_reg, col_reg}<22'b0110110000101101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b0110110000101101111110) && ({row_reg, col_reg}<22'b0110110000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110000110000000010) && ({row_reg, col_reg}<22'b0110110000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110000110000101101) && ({row_reg, col_reg}<22'b0110110001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110001000001010111) && ({row_reg, col_reg}<22'b0110110001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110001000010000010) && ({row_reg, col_reg}<22'b0110110001000100000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110001000100000110) && ({row_reg, col_reg}<22'b0110110001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110001001000000010) && ({row_reg, col_reg}<22'b0110110001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110001001010000010) && ({row_reg, col_reg}<22'b0110110001001101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001001101111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110001001101111110) && ({row_reg, col_reg}<22'b0110110001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110001010000000010) && ({row_reg, col_reg}<22'b0110110001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110001010000101101) && ({row_reg, col_reg}<22'b0110110001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110001100001010111) && ({row_reg, col_reg}<22'b0110110001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110001100010000010) && ({row_reg, col_reg}<22'b0110110001100100000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110001100100000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110110001100100000111) && ({row_reg, col_reg}<22'b0110110001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110001101000000010) && ({row_reg, col_reg}<22'b0110110001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110001101010000010) && ({row_reg, col_reg}<22'b0110110001101101111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001101101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110110001101101111101) && ({row_reg, col_reg}<22'b0110110001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110001110000000010) && ({row_reg, col_reg}<22'b0110110001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110001110000101101) && ({row_reg, col_reg}<22'b0110110010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110010000001010111) && ({row_reg, col_reg}<22'b0110110010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110010000010000010) && ({row_reg, col_reg}<22'b0110110010000100000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110010000100000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110010000100001000) && ({row_reg, col_reg}<22'b0110110010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110010001000000010) && ({row_reg, col_reg}<22'b0110110010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110010001010000010) && ({row_reg, col_reg}<22'b0110110010001101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010001101111011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b0110110010001101111100) && ({row_reg, col_reg}<22'b0110110010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110010010000000010) && ({row_reg, col_reg}<22'b0110110010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110010010000101101) && ({row_reg, col_reg}<22'b0110110010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110010100001010111) && ({row_reg, col_reg}<22'b0110110010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110010100010000010) && ({row_reg, col_reg}<22'b0110110010100100001000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110010100100001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110010100100001001) && ({row_reg, col_reg}<22'b0110110010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110010101000000010) && ({row_reg, col_reg}<22'b0110110010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110010101010000010) && ({row_reg, col_reg}<22'b0110110010101101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010101101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110110010101101111011) && ({row_reg, col_reg}<22'b0110110010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110010110000000010) && ({row_reg, col_reg}<22'b0110110010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110010110000101101) && ({row_reg, col_reg}<22'b0110110011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110011000001010111) && ({row_reg, col_reg}<22'b0110110011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110011000010000010) && ({row_reg, col_reg}<22'b0110110011000100001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110011000100001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110110011000100001010) && ({row_reg, col_reg}<22'b0110110011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110011001000000010) && ({row_reg, col_reg}<22'b0110110011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110011001010000010) && ({row_reg, col_reg}<22'b0110110011001101111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011001101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0110110011001101111010) && ({row_reg, col_reg}<22'b0110110011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110011010000000010) && ({row_reg, col_reg}<22'b0110110011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110011010000101101) && ({row_reg, col_reg}<22'b0110110011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110011100001010111) && ({row_reg, col_reg}<22'b0110110011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110011100010000010) && ({row_reg, col_reg}<22'b0110110011100100001011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110011100100001011) && ({row_reg, col_reg}<22'b0110110011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110011101000000010) && ({row_reg, col_reg}<22'b0110110011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110011101010000010) && ({row_reg, col_reg}<22'b0110110011101101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011101101111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110110011101101111001) && ({row_reg, col_reg}<22'b0110110011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110011110000000010) && ({row_reg, col_reg}<22'b0110110011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110011110000101101) && ({row_reg, col_reg}<22'b0110110100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110100000001010111) && ({row_reg, col_reg}<22'b0110110100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110100000010000010) && ({row_reg, col_reg}<22'b0110110100000100001100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110100000100001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110110100000100001101) && ({row_reg, col_reg}<22'b0110110100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110110100001000000010) && ({row_reg, col_reg}<22'b0110110100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110100001010000010) && ({row_reg, col_reg}<22'b0110110100001101110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100001101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0110110100001101110111) && ({row_reg, col_reg}<22'b0110110100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110100010000000010) && ({row_reg, col_reg}<22'b0110110100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110100010000101101) && ({row_reg, col_reg}<22'b0110110100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110100100001010111) && ({row_reg, col_reg}<22'b0110110100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110100100010000010) && ({row_reg, col_reg}<22'b0110110100100100001110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110100100100001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110110100100100001111) && ({row_reg, col_reg}<22'b0110110100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110110100101000000010) && ({row_reg, col_reg}<22'b0110110100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110100101010000010) && ({row_reg, col_reg}<22'b0110110100101101110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100101101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b0110110100101101110101) && ({row_reg, col_reg}<22'b0110110100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110100110000000010) && ({row_reg, col_reg}<22'b0110110100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110100110000101101) && ({row_reg, col_reg}<22'b0110110101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110101000001010111) && ({row_reg, col_reg}<22'b0110110101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110101000010000010) && ({row_reg, col_reg}<22'b0110110101000100010000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110101000100010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==22'b0110110101000100010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b0110110101000100010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0110110101000100010011) && ({row_reg, col_reg}<22'b0110110101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110110101001000000010) && ({row_reg, col_reg}<22'b0110110101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110101001010000010) && ({row_reg, col_reg}<22'b0110110101001101110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101001101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b0110110101001101110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b0110110101001101110011) && ({row_reg, col_reg}<22'b0110110101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110101010000000010) && ({row_reg, col_reg}<22'b0110110101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110101010000101101) && ({row_reg, col_reg}<22'b0110110101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110101100001010111) && ({row_reg, col_reg}<22'b0110110101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110101100010000010) && ({row_reg, col_reg}<22'b0110110101100100010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110101100100010110) && ({row_reg, col_reg}<22'b0110110101100111010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110101100111010111) && ({row_reg, col_reg}<22'b0110110101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110110101101000000010) && ({row_reg, col_reg}<22'b0110110101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110101101010000010) && ({row_reg, col_reg}<22'b0110110101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101101010101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b0110110101101010101101) && ({row_reg, col_reg}<22'b0110110101101101101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110101101101101101) && ({row_reg, col_reg}<22'b0110110101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110101110000000010) && ({row_reg, col_reg}<22'b0110110101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110101110000101101) && ({row_reg, col_reg}<22'b0110110110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110110000001010111) && ({row_reg, col_reg}<22'b0110110110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110110110000010000010) && ({row_reg, col_reg}<22'b0110110110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110110000111010111) && ({row_reg, col_reg}<22'b0110110110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110110110001000000010) && ({row_reg, col_reg}<22'b0110110110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110110001010000010) && ({row_reg, col_reg}<22'b0110110110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110110001010101101) && ({row_reg, col_reg}<22'b0110110110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110110010000000010) && ({row_reg, col_reg}<22'b0110110110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110110010000101101) && ({row_reg, col_reg}<22'b0110110110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110110100001010111) && ({row_reg, col_reg}<22'b0110110110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110110110100010000010) && ({row_reg, col_reg}<22'b0110110110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110110100111010111) && ({row_reg, col_reg}<22'b0110110110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110110110101000000010) && ({row_reg, col_reg}<22'b0110110110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110110101010000010) && ({row_reg, col_reg}<22'b0110110110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110110101010101101) && ({row_reg, col_reg}<22'b0110110110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110110110000000010) && ({row_reg, col_reg}<22'b0110110110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110110110000101101) && ({row_reg, col_reg}<22'b0110110111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110111000001010111) && ({row_reg, col_reg}<22'b0110110111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110110111000010000010) && ({row_reg, col_reg}<22'b0110110111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110111000111010111) && ({row_reg, col_reg}<22'b0110110111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110110111001000000010) && ({row_reg, col_reg}<22'b0110110111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110111001010000010) && ({row_reg, col_reg}<22'b0110110111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110111001010101101) && ({row_reg, col_reg}<22'b0110110111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110111010000000010) && ({row_reg, col_reg}<22'b0110110111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110111010000101101) && ({row_reg, col_reg}<22'b0110110111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110111100001010111) && ({row_reg, col_reg}<22'b0110110111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110110111100010000010) && ({row_reg, col_reg}<22'b0110110111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110110111100111010111) && ({row_reg, col_reg}<22'b0110110111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110110111101000000010) && ({row_reg, col_reg}<22'b0110110111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110111101010000010) && ({row_reg, col_reg}<22'b0110110111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110111101010101101) && ({row_reg, col_reg}<22'b0110110111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110110111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110110111110000000010) && ({row_reg, col_reg}<22'b0110110111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110110111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110110111110000101101) && ({row_reg, col_reg}<22'b0110111000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111000000001010111) && ({row_reg, col_reg}<22'b0110111000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110111000000010000010) && ({row_reg, col_reg}<22'b0110111000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111000000111010111) && ({row_reg, col_reg}<22'b0110111000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111000001000000010) && ({row_reg, col_reg}<22'b0110111000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111000001010000010) && ({row_reg, col_reg}<22'b0110111000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111000001010101101) && ({row_reg, col_reg}<22'b0110111000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111000010000000010) && ({row_reg, col_reg}<22'b0110111000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111000010000101101) && ({row_reg, col_reg}<22'b0110111000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111000100001010111) && ({row_reg, col_reg}<22'b0110111000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110111000100010000010) && ({row_reg, col_reg}<22'b0110111000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111000100111010111) && ({row_reg, col_reg}<22'b0110111000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111000101000000010) && ({row_reg, col_reg}<22'b0110111000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111000101010000010) && ({row_reg, col_reg}<22'b0110111000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111000101010101101) && ({row_reg, col_reg}<22'b0110111000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111000110000000010) && ({row_reg, col_reg}<22'b0110111000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111000110000101101) && ({row_reg, col_reg}<22'b0110111001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111001000001010111) && ({row_reg, col_reg}<22'b0110111001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110111001000010000010) && ({row_reg, col_reg}<22'b0110111001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111001000111010111) && ({row_reg, col_reg}<22'b0110111001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111001001000000010) && ({row_reg, col_reg}<22'b0110111001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111001001010000010) && ({row_reg, col_reg}<22'b0110111001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111001001010101101) && ({row_reg, col_reg}<22'b0110111001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111001010000000010) && ({row_reg, col_reg}<22'b0110111001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111001010000101101) && ({row_reg, col_reg}<22'b0110111001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111001100001010111) && ({row_reg, col_reg}<22'b0110111001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111001100010000010) && ({row_reg, col_reg}<22'b0110111001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111001100111010111) && ({row_reg, col_reg}<22'b0110111001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111001101000000010) && ({row_reg, col_reg}<22'b0110111001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111001101010000010) && ({row_reg, col_reg}<22'b0110111001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111001101010101101) && ({row_reg, col_reg}<22'b0110111001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111001110000000010) && ({row_reg, col_reg}<22'b0110111001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111001110000101101) && ({row_reg, col_reg}<22'b0110111010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111010000001010111) && ({row_reg, col_reg}<22'b0110111010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111010000010000010) && ({row_reg, col_reg}<22'b0110111010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111010000111010111) && ({row_reg, col_reg}<22'b0110111010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111010001000000010) && ({row_reg, col_reg}<22'b0110111010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111010001010000010) && ({row_reg, col_reg}<22'b0110111010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111010001010101101) && ({row_reg, col_reg}<22'b0110111010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111010010000000010) && ({row_reg, col_reg}<22'b0110111010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111010010000101101) && ({row_reg, col_reg}<22'b0110111010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111010100001010111) && ({row_reg, col_reg}<22'b0110111010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111010100010000010) && ({row_reg, col_reg}<22'b0110111010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111010100111010111) && ({row_reg, col_reg}<22'b0110111010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111010101000000010) && ({row_reg, col_reg}<22'b0110111010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111010101010000010) && ({row_reg, col_reg}<22'b0110111010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111010101010101101) && ({row_reg, col_reg}<22'b0110111010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111010110000000010) && ({row_reg, col_reg}<22'b0110111010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111010110000101101) && ({row_reg, col_reg}<22'b0110111011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111011000001010111) && ({row_reg, col_reg}<22'b0110111011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111011000010000010) && ({row_reg, col_reg}<22'b0110111011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111011000111010111) && ({row_reg, col_reg}<22'b0110111011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111011001000000010) && ({row_reg, col_reg}<22'b0110111011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111011001010000010) && ({row_reg, col_reg}<22'b0110111011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111011001010101101) && ({row_reg, col_reg}<22'b0110111011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111011010000000010) && ({row_reg, col_reg}<22'b0110111011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111011010000101101) && ({row_reg, col_reg}<22'b0110111011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111011100001010111) && ({row_reg, col_reg}<22'b0110111011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111011100010000010) && ({row_reg, col_reg}<22'b0110111011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111011100111010111) && ({row_reg, col_reg}<22'b0110111011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111011101000000010) && ({row_reg, col_reg}<22'b0110111011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111011101010000010) && ({row_reg, col_reg}<22'b0110111011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111011101010101101) && ({row_reg, col_reg}<22'b0110111011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111011110000000010) && ({row_reg, col_reg}<22'b0110111011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111011110000101101) && ({row_reg, col_reg}<22'b0110111100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111100000001010111) && ({row_reg, col_reg}<22'b0110111100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111100000010000010) && ({row_reg, col_reg}<22'b0110111100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111100000111010111) && ({row_reg, col_reg}<22'b0110111100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111100001000000010) && ({row_reg, col_reg}<22'b0110111100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111100001010000010) && ({row_reg, col_reg}<22'b0110111100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111100001010101101) && ({row_reg, col_reg}<22'b0110111100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111100010000000010) && ({row_reg, col_reg}<22'b0110111100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111100010000101101) && ({row_reg, col_reg}<22'b0110111100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111100100001010111) && ({row_reg, col_reg}<22'b0110111100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111100100010000010) && ({row_reg, col_reg}<22'b0110111100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111100100111010111) && ({row_reg, col_reg}<22'b0110111100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111100101000000010) && ({row_reg, col_reg}<22'b0110111100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111100101010000010) && ({row_reg, col_reg}<22'b0110111100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111100101010101101) && ({row_reg, col_reg}<22'b0110111100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111100110000000010) && ({row_reg, col_reg}<22'b0110111100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111100110000101101) && ({row_reg, col_reg}<22'b0110111101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111101000001010111) && ({row_reg, col_reg}<22'b0110111101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111101000010000010) && ({row_reg, col_reg}<22'b0110111101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111101000111010111) && ({row_reg, col_reg}<22'b0110111101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111101001000000010) && ({row_reg, col_reg}<22'b0110111101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111101001010000010) && ({row_reg, col_reg}<22'b0110111101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111101001010101101) && ({row_reg, col_reg}<22'b0110111101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111101010000000010) && ({row_reg, col_reg}<22'b0110111101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111101010000101101) && ({row_reg, col_reg}<22'b0110111101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111101100001010111) && ({row_reg, col_reg}<22'b0110111101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111101100010000010) && ({row_reg, col_reg}<22'b0110111101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111101100111010111) && ({row_reg, col_reg}<22'b0110111101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111101101000000010) && ({row_reg, col_reg}<22'b0110111101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111101101010000010) && ({row_reg, col_reg}<22'b0110111101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111101101010101101) && ({row_reg, col_reg}<22'b0110111101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111101110000000010) && ({row_reg, col_reg}<22'b0110111101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111101110000101101) && ({row_reg, col_reg}<22'b0110111110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111110000001010111) && ({row_reg, col_reg}<22'b0110111110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111110000010000010) && ({row_reg, col_reg}<22'b0110111110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111110000111010111) && ({row_reg, col_reg}<22'b0110111110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110111110001000000010) && ({row_reg, col_reg}<22'b0110111110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111110001010000010) && ({row_reg, col_reg}<22'b0110111110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111110001010101101) && ({row_reg, col_reg}<22'b0110111110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111110010000000010) && ({row_reg, col_reg}<22'b0110111110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111110010000101101) && ({row_reg, col_reg}<22'b0110111110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111110100001010111) && ({row_reg, col_reg}<22'b0110111110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111110100010000010) && ({row_reg, col_reg}<22'b0110111110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111110100111010111) && ({row_reg, col_reg}<22'b0110111110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0110111110101000000010) && ({row_reg, col_reg}<22'b0110111110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111110101010000010) && ({row_reg, col_reg}<22'b0110111110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111110101010101101) && ({row_reg, col_reg}<22'b0110111110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111110110000000010) && ({row_reg, col_reg}<22'b0110111110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111110110000101101) && ({row_reg, col_reg}<22'b0110111111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111111000001010111) && ({row_reg, col_reg}<22'b0110111111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111111000010000010) && ({row_reg, col_reg}<22'b0110111111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111111000111010111) && ({row_reg, col_reg}<22'b0110111111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110111111001000000010) && ({row_reg, col_reg}<22'b0110111111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111111001010000010) && ({row_reg, col_reg}<22'b0110111111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111111001010101101) && ({row_reg, col_reg}<22'b0110111111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111111010000000010) && ({row_reg, col_reg}<22'b0110111111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111111010000101101) && ({row_reg, col_reg}<22'b0110111111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111111100001010111) && ({row_reg, col_reg}<22'b0110111111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0110111111100010000010) && ({row_reg, col_reg}<22'b0110111111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0110111111100111010111) && ({row_reg, col_reg}<22'b0110111111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0110111111101000000010) && ({row_reg, col_reg}<22'b0110111111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111111101010000010) && ({row_reg, col_reg}<22'b0110111111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111111101010101101) && ({row_reg, col_reg}<22'b0110111111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0110111111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0110111111110000000010) && ({row_reg, col_reg}<22'b0110111111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0110111111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0110111111110000101101) && ({row_reg, col_reg}<22'b0111000000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000000000001010111) && ({row_reg, col_reg}<22'b0111000000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111000000000010000010) && ({row_reg, col_reg}<22'b0111000000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000000000111010111) && ({row_reg, col_reg}<22'b0111000000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111000000001000000010) && ({row_reg, col_reg}<22'b0111000000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000000001010000010) && ({row_reg, col_reg}<22'b0111000000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000000001010101101) && ({row_reg, col_reg}<22'b0111000000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000000010000000010) && ({row_reg, col_reg}<22'b0111000000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000000010000101101) && ({row_reg, col_reg}<22'b0111000000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000000100001010111) && ({row_reg, col_reg}<22'b0111000000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111000000100010000010) && ({row_reg, col_reg}<22'b0111000000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000000100111010111) && ({row_reg, col_reg}<22'b0111000000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111000000101000000010) && ({row_reg, col_reg}<22'b0111000000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000000101010000010) && ({row_reg, col_reg}<22'b0111000000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000000101010101101) && ({row_reg, col_reg}<22'b0111000000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000000110000000010) && ({row_reg, col_reg}<22'b0111000000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000000110000101101) && ({row_reg, col_reg}<22'b0111000001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000001000001010111) && ({row_reg, col_reg}<22'b0111000001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111000001000010000010) && ({row_reg, col_reg}<22'b0111000001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000001000111010111) && ({row_reg, col_reg}<22'b0111000001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111000001001000000010) && ({row_reg, col_reg}<22'b0111000001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000001001010000010) && ({row_reg, col_reg}<22'b0111000001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000001001010101101) && ({row_reg, col_reg}<22'b0111000001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000001010000000010) && ({row_reg, col_reg}<22'b0111000001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000001010000101101) && ({row_reg, col_reg}<22'b0111000001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000001100001010111) && ({row_reg, col_reg}<22'b0111000001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111000001100010000010) && ({row_reg, col_reg}<22'b0111000001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000001100111010111) && ({row_reg, col_reg}<22'b0111000001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000001101000000010) && ({row_reg, col_reg}<22'b0111000001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000001101010000010) && ({row_reg, col_reg}<22'b0111000001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000001101010101101) && ({row_reg, col_reg}<22'b0111000001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000001110000000010) && ({row_reg, col_reg}<22'b0111000001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000001110000101101) && ({row_reg, col_reg}<22'b0111000010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000010000001010111) && ({row_reg, col_reg}<22'b0111000010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111000010000010000010) && ({row_reg, col_reg}<22'b0111000010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000010000111010111) && ({row_reg, col_reg}<22'b0111000010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000010001000000010) && ({row_reg, col_reg}<22'b0111000010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000010001010000010) && ({row_reg, col_reg}<22'b0111000010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000010001010101101) && ({row_reg, col_reg}<22'b0111000010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000010010000000010) && ({row_reg, col_reg}<22'b0111000010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000010010000101101) && ({row_reg, col_reg}<22'b0111000010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000010100001010111) && ({row_reg, col_reg}<22'b0111000010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111000010100010000010) && ({row_reg, col_reg}<22'b0111000010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000010100111010111) && ({row_reg, col_reg}<22'b0111000010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000010101000000010) && ({row_reg, col_reg}<22'b0111000010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000010101010000010) && ({row_reg, col_reg}<22'b0111000010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000010101010101101) && ({row_reg, col_reg}<22'b0111000010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000010110000000010) && ({row_reg, col_reg}<22'b0111000010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000010110000101101) && ({row_reg, col_reg}<22'b0111000011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000011000001010111) && ({row_reg, col_reg}<22'b0111000011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111000011000010000010) && ({row_reg, col_reg}<22'b0111000011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000011000111010111) && ({row_reg, col_reg}<22'b0111000011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000011001000000010) && ({row_reg, col_reg}<22'b0111000011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000011001010000010) && ({row_reg, col_reg}<22'b0111000011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000011001010101101) && ({row_reg, col_reg}<22'b0111000011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000011010000000010) && ({row_reg, col_reg}<22'b0111000011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000011010000101101) && ({row_reg, col_reg}<22'b0111000011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000011100001010111) && ({row_reg, col_reg}<22'b0111000011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000011100010000010) && ({row_reg, col_reg}<22'b0111000011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000011100111010111) && ({row_reg, col_reg}<22'b0111000011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000011101000000010) && ({row_reg, col_reg}<22'b0111000011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000011101010000010) && ({row_reg, col_reg}<22'b0111000011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000011101010101101) && ({row_reg, col_reg}<22'b0111000011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000011110000000010) && ({row_reg, col_reg}<22'b0111000011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000011110000101101) && ({row_reg, col_reg}<22'b0111000100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000100000001010111) && ({row_reg, col_reg}<22'b0111000100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000100000010000010) && ({row_reg, col_reg}<22'b0111000100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000100000111010111) && ({row_reg, col_reg}<22'b0111000100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000100001000000010) && ({row_reg, col_reg}<22'b0111000100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000100001010000010) && ({row_reg, col_reg}<22'b0111000100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000100001010101101) && ({row_reg, col_reg}<22'b0111000100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000100010000000010) && ({row_reg, col_reg}<22'b0111000100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000100010000101101) && ({row_reg, col_reg}<22'b0111000100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000100100001010111) && ({row_reg, col_reg}<22'b0111000100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000100100010000010) && ({row_reg, col_reg}<22'b0111000100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000100100111010111) && ({row_reg, col_reg}<22'b0111000100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000100101000000010) && ({row_reg, col_reg}<22'b0111000100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000100101010000010) && ({row_reg, col_reg}<22'b0111000100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000100101010101101) && ({row_reg, col_reg}<22'b0111000100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000100110000000010) && ({row_reg, col_reg}<22'b0111000100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000100110000101101) && ({row_reg, col_reg}<22'b0111000101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000101000001010111) && ({row_reg, col_reg}<22'b0111000101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000101000010000010) && ({row_reg, col_reg}<22'b0111000101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000101000111010111) && ({row_reg, col_reg}<22'b0111000101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000101001000000010) && ({row_reg, col_reg}<22'b0111000101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000101001010000010) && ({row_reg, col_reg}<22'b0111000101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000101001010101101) && ({row_reg, col_reg}<22'b0111000101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000101010000000010) && ({row_reg, col_reg}<22'b0111000101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000101010000101101) && ({row_reg, col_reg}<22'b0111000101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000101100001010111) && ({row_reg, col_reg}<22'b0111000101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000101100010000010) && ({row_reg, col_reg}<22'b0111000101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000101100111010111) && ({row_reg, col_reg}<22'b0111000101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000101101000000010) && ({row_reg, col_reg}<22'b0111000101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000101101010000010) && ({row_reg, col_reg}<22'b0111000101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000101101010101101) && ({row_reg, col_reg}<22'b0111000101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000101110000000010) && ({row_reg, col_reg}<22'b0111000101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000101110000101101) && ({row_reg, col_reg}<22'b0111000110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000110000001010111) && ({row_reg, col_reg}<22'b0111000110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000110000010000010) && ({row_reg, col_reg}<22'b0111000110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000110000111010111) && ({row_reg, col_reg}<22'b0111000110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000110001000000010) && ({row_reg, col_reg}<22'b0111000110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000110001010000010) && ({row_reg, col_reg}<22'b0111000110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000110001010101101) && ({row_reg, col_reg}<22'b0111000110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000110010000000010) && ({row_reg, col_reg}<22'b0111000110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000110010000101101) && ({row_reg, col_reg}<22'b0111000110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000110100001010111) && ({row_reg, col_reg}<22'b0111000110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000110100010000010) && ({row_reg, col_reg}<22'b0111000110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000110100111010111) && ({row_reg, col_reg}<22'b0111000110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000110101000000010) && ({row_reg, col_reg}<22'b0111000110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000110101010000010) && ({row_reg, col_reg}<22'b0111000110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000110101010101101) && ({row_reg, col_reg}<22'b0111000110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000110110000000010) && ({row_reg, col_reg}<22'b0111000110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000110110000101101) && ({row_reg, col_reg}<22'b0111000111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000111000001010111) && ({row_reg, col_reg}<22'b0111000111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000111000010000010) && ({row_reg, col_reg}<22'b0111000111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000111000111010111) && ({row_reg, col_reg}<22'b0111000111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000111001000000010) && ({row_reg, col_reg}<22'b0111000111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000111001010000010) && ({row_reg, col_reg}<22'b0111000111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000111001010101101) && ({row_reg, col_reg}<22'b0111000111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000111010000000010) && ({row_reg, col_reg}<22'b0111000111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000111010000101101) && ({row_reg, col_reg}<22'b0111000111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000111100001010111) && ({row_reg, col_reg}<22'b0111000111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000111100010000010) && ({row_reg, col_reg}<22'b0111000111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111000111100111010111) && ({row_reg, col_reg}<22'b0111000111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111000111101000000010) && ({row_reg, col_reg}<22'b0111000111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000111101010000010) && ({row_reg, col_reg}<22'b0111000111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000111101010101101) && ({row_reg, col_reg}<22'b0111000111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111000111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111000111110000000010) && ({row_reg, col_reg}<22'b0111000111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111000111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111000111110000101101) && ({row_reg, col_reg}<22'b0111001000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001000000001010111) && ({row_reg, col_reg}<22'b0111001000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001000000010000010) && ({row_reg, col_reg}<22'b0111001000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001000000111010111) && ({row_reg, col_reg}<22'b0111001000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001000001000000010) && ({row_reg, col_reg}<22'b0111001000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001000001010000010) && ({row_reg, col_reg}<22'b0111001000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001000001010101101) && ({row_reg, col_reg}<22'b0111001000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001000010000000010) && ({row_reg, col_reg}<22'b0111001000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001000010000101101) && ({row_reg, col_reg}<22'b0111001000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001000100001010111) && ({row_reg, col_reg}<22'b0111001000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001000100010000010) && ({row_reg, col_reg}<22'b0111001000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001000100111010111) && ({row_reg, col_reg}<22'b0111001000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001000101000000010) && ({row_reg, col_reg}<22'b0111001000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001000101010000010) && ({row_reg, col_reg}<22'b0111001000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001000101010101101) && ({row_reg, col_reg}<22'b0111001000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001000110000000010) && ({row_reg, col_reg}<22'b0111001000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001000110000101101) && ({row_reg, col_reg}<22'b0111001001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001001000001010111) && ({row_reg, col_reg}<22'b0111001001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001001000010000010) && ({row_reg, col_reg}<22'b0111001001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001001000111010111) && ({row_reg, col_reg}<22'b0111001001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111001001001000000010) && ({row_reg, col_reg}<22'b0111001001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001001001010000010) && ({row_reg, col_reg}<22'b0111001001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001001001010101101) && ({row_reg, col_reg}<22'b0111001001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001001010000000010) && ({row_reg, col_reg}<22'b0111001001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001001010000101101) && ({row_reg, col_reg}<22'b0111001001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001001100001010111) && ({row_reg, col_reg}<22'b0111001001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001001100010000010) && ({row_reg, col_reg}<22'b0111001001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001001100111010111) && ({row_reg, col_reg}<22'b0111001001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111001001101000000010) && ({row_reg, col_reg}<22'b0111001001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001001101010000010) && ({row_reg, col_reg}<22'b0111001001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001001101010101101) && ({row_reg, col_reg}<22'b0111001001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001001110000000010) && ({row_reg, col_reg}<22'b0111001001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001001110000101101) && ({row_reg, col_reg}<22'b0111001010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001010000001010111) && ({row_reg, col_reg}<22'b0111001010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001010000010000010) && ({row_reg, col_reg}<22'b0111001010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001010000111010111) && ({row_reg, col_reg}<22'b0111001010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111001010001000000010) && ({row_reg, col_reg}<22'b0111001010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001010001010000010) && ({row_reg, col_reg}<22'b0111001010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001010001010101101) && ({row_reg, col_reg}<22'b0111001010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001010010000000010) && ({row_reg, col_reg}<22'b0111001010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001010010000101101) && ({row_reg, col_reg}<22'b0111001010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001010100001010111) && ({row_reg, col_reg}<22'b0111001010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001010100010000010) && ({row_reg, col_reg}<22'b0111001010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001010100111010111) && ({row_reg, col_reg}<22'b0111001010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001010101000000010) && ({row_reg, col_reg}<22'b0111001010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001010101010000010) && ({row_reg, col_reg}<22'b0111001010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001010101010101101) && ({row_reg, col_reg}<22'b0111001010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001010110000000010) && ({row_reg, col_reg}<22'b0111001010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001010110000101101) && ({row_reg, col_reg}<22'b0111001011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001011000001010111) && ({row_reg, col_reg}<22'b0111001011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111001011000010000010) && ({row_reg, col_reg}<22'b0111001011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001011000111010111) && ({row_reg, col_reg}<22'b0111001011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001011001000000010) && ({row_reg, col_reg}<22'b0111001011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001011001010000010) && ({row_reg, col_reg}<22'b0111001011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001011001010101101) && ({row_reg, col_reg}<22'b0111001011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001011010000000010) && ({row_reg, col_reg}<22'b0111001011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001011010000101101) && ({row_reg, col_reg}<22'b0111001011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001011100001010111) && ({row_reg, col_reg}<22'b0111001011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111001011100010000010) && ({row_reg, col_reg}<22'b0111001011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001011100111010111) && ({row_reg, col_reg}<22'b0111001011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001011101000000010) && ({row_reg, col_reg}<22'b0111001011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001011101010000010) && ({row_reg, col_reg}<22'b0111001011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001011101010101101) && ({row_reg, col_reg}<22'b0111001011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001011110000000010) && ({row_reg, col_reg}<22'b0111001011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001011110000101101) && ({row_reg, col_reg}<22'b0111001100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001100000001010111) && ({row_reg, col_reg}<22'b0111001100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111001100000010000010) && ({row_reg, col_reg}<22'b0111001100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001100000111010111) && ({row_reg, col_reg}<22'b0111001100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001100001000000010) && ({row_reg, col_reg}<22'b0111001100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001100001010000010) && ({row_reg, col_reg}<22'b0111001100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001100001010101101) && ({row_reg, col_reg}<22'b0111001100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001100010000000010) && ({row_reg, col_reg}<22'b0111001100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001100010000101101) && ({row_reg, col_reg}<22'b0111001100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001100100001010111) && ({row_reg, col_reg}<22'b0111001100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001100100010000010) && ({row_reg, col_reg}<22'b0111001100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001100100111010111) && ({row_reg, col_reg}<22'b0111001100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001100101000000010) && ({row_reg, col_reg}<22'b0111001100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001100101010000010) && ({row_reg, col_reg}<22'b0111001100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001100101010101101) && ({row_reg, col_reg}<22'b0111001100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001100110000000010) && ({row_reg, col_reg}<22'b0111001100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001100110000101101) && ({row_reg, col_reg}<22'b0111001101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001101000001010111) && ({row_reg, col_reg}<22'b0111001101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111001101000010000010) && ({row_reg, col_reg}<22'b0111001101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001101000111010111) && ({row_reg, col_reg}<22'b0111001101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001101001000000010) && ({row_reg, col_reg}<22'b0111001101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001101001010000010) && ({row_reg, col_reg}<22'b0111001101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001101001010101101) && ({row_reg, col_reg}<22'b0111001101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001101010000000010) && ({row_reg, col_reg}<22'b0111001101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001101010000101101) && ({row_reg, col_reg}<22'b0111001101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001101100001010111) && ({row_reg, col_reg}<22'b0111001101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001101100010000010) && ({row_reg, col_reg}<22'b0111001101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001101100111010111) && ({row_reg, col_reg}<22'b0111001101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001101101000000010) && ({row_reg, col_reg}<22'b0111001101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001101101010000010) && ({row_reg, col_reg}<22'b0111001101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001101101010101101) && ({row_reg, col_reg}<22'b0111001101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001101110000000010) && ({row_reg, col_reg}<22'b0111001101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001101110000101101) && ({row_reg, col_reg}<22'b0111001110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001110000001010111) && ({row_reg, col_reg}<22'b0111001110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001110000010000010) && ({row_reg, col_reg}<22'b0111001110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001110000111010111) && ({row_reg, col_reg}<22'b0111001110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001110001000000010) && ({row_reg, col_reg}<22'b0111001110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001110001010000010) && ({row_reg, col_reg}<22'b0111001110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001110001010101101) && ({row_reg, col_reg}<22'b0111001110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001110010000000010) && ({row_reg, col_reg}<22'b0111001110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001110010000101101) && ({row_reg, col_reg}<22'b0111001110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001110100001010111) && ({row_reg, col_reg}<22'b0111001110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001110100010000010) && ({row_reg, col_reg}<22'b0111001110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001110100111010111) && ({row_reg, col_reg}<22'b0111001110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001110101000000010) && ({row_reg, col_reg}<22'b0111001110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001110101010000010) && ({row_reg, col_reg}<22'b0111001110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001110101010101101) && ({row_reg, col_reg}<22'b0111001110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001110110000000010) && ({row_reg, col_reg}<22'b0111001110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001110110000101101) && ({row_reg, col_reg}<22'b0111001111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001111000001010111) && ({row_reg, col_reg}<22'b0111001111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001111000010000010) && ({row_reg, col_reg}<22'b0111001111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001111000111010111) && ({row_reg, col_reg}<22'b0111001111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001111001000000010) && ({row_reg, col_reg}<22'b0111001111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001111001010000010) && ({row_reg, col_reg}<22'b0111001111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001111001010101101) && ({row_reg, col_reg}<22'b0111001111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001111010000000010) && ({row_reg, col_reg}<22'b0111001111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001111010000101101) && ({row_reg, col_reg}<22'b0111001111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001111100001010111) && ({row_reg, col_reg}<22'b0111001111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001111100010000010) && ({row_reg, col_reg}<22'b0111001111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111001111100111010111) && ({row_reg, col_reg}<22'b0111001111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111001111101000000010) && ({row_reg, col_reg}<22'b0111001111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001111101010000010) && ({row_reg, col_reg}<22'b0111001111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001111101010101101) && ({row_reg, col_reg}<22'b0111001111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111001111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111001111110000000010) && ({row_reg, col_reg}<22'b0111001111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111001111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111001111110000101101) && ({row_reg, col_reg}<22'b0111010000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010000000001010111) && ({row_reg, col_reg}<22'b0111010000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010000000010000010) && ({row_reg, col_reg}<22'b0111010000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010000000111010111) && ({row_reg, col_reg}<22'b0111010000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010000001000000010) && ({row_reg, col_reg}<22'b0111010000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010000001010000010) && ({row_reg, col_reg}<22'b0111010000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010000001010101101) && ({row_reg, col_reg}<22'b0111010000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010000010000000010) && ({row_reg, col_reg}<22'b0111010000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010000010000101101) && ({row_reg, col_reg}<22'b0111010000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010000100001010111) && ({row_reg, col_reg}<22'b0111010000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010000100010000010) && ({row_reg, col_reg}<22'b0111010000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010000100111010111) && ({row_reg, col_reg}<22'b0111010000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010000101000000010) && ({row_reg, col_reg}<22'b0111010000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010000101010000010) && ({row_reg, col_reg}<22'b0111010000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010000101010101101) && ({row_reg, col_reg}<22'b0111010000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010000110000000010) && ({row_reg, col_reg}<22'b0111010000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010000110000101101) && ({row_reg, col_reg}<22'b0111010001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010001000001010111) && ({row_reg, col_reg}<22'b0111010001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010001000010000010) && ({row_reg, col_reg}<22'b0111010001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010001000111010111) && ({row_reg, col_reg}<22'b0111010001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010001001000000010) && ({row_reg, col_reg}<22'b0111010001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010001001010000010) && ({row_reg, col_reg}<22'b0111010001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010001001010101101) && ({row_reg, col_reg}<22'b0111010001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010001010000000010) && ({row_reg, col_reg}<22'b0111010001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010001010000101101) && ({row_reg, col_reg}<22'b0111010001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010001100001010111) && ({row_reg, col_reg}<22'b0111010001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010001100010000010) && ({row_reg, col_reg}<22'b0111010001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010001100111010111) && ({row_reg, col_reg}<22'b0111010001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010001101000000010) && ({row_reg, col_reg}<22'b0111010001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010001101010000010) && ({row_reg, col_reg}<22'b0111010001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010001101010101101) && ({row_reg, col_reg}<22'b0111010001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010001110000000010) && ({row_reg, col_reg}<22'b0111010001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010001110000101101) && ({row_reg, col_reg}<22'b0111010010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010010000001010111) && ({row_reg, col_reg}<22'b0111010010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010010000010000010) && ({row_reg, col_reg}<22'b0111010010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010010000111010111) && ({row_reg, col_reg}<22'b0111010010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010010001000000010) && ({row_reg, col_reg}<22'b0111010010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010010001010000010) && ({row_reg, col_reg}<22'b0111010010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010010001010101101) && ({row_reg, col_reg}<22'b0111010010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010010010000000010) && ({row_reg, col_reg}<22'b0111010010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010010010000101101) && ({row_reg, col_reg}<22'b0111010010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010010100001010111) && ({row_reg, col_reg}<22'b0111010010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010010100010000010) && ({row_reg, col_reg}<22'b0111010010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010010100111010111) && ({row_reg, col_reg}<22'b0111010010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010010101000000010) && ({row_reg, col_reg}<22'b0111010010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010010101010000010) && ({row_reg, col_reg}<22'b0111010010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010010101010101101) && ({row_reg, col_reg}<22'b0111010010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010010110000000010) && ({row_reg, col_reg}<22'b0111010010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010010110000101101) && ({row_reg, col_reg}<22'b0111010011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010011000001010111) && ({row_reg, col_reg}<22'b0111010011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010011000010000010) && ({row_reg, col_reg}<22'b0111010011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010011000111010111) && ({row_reg, col_reg}<22'b0111010011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111010011001000000010) && ({row_reg, col_reg}<22'b0111010011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010011001010000010) && ({row_reg, col_reg}<22'b0111010011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010011001010101101) && ({row_reg, col_reg}<22'b0111010011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010011010000000010) && ({row_reg, col_reg}<22'b0111010011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010011010000101101) && ({row_reg, col_reg}<22'b0111010011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010011100001010111) && ({row_reg, col_reg}<22'b0111010011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010011100010000010) && ({row_reg, col_reg}<22'b0111010011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010011100111010111) && ({row_reg, col_reg}<22'b0111010011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111010011101000000010) && ({row_reg, col_reg}<22'b0111010011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010011101010000010) && ({row_reg, col_reg}<22'b0111010011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010011101010101101) && ({row_reg, col_reg}<22'b0111010011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010011110000000010) && ({row_reg, col_reg}<22'b0111010011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010011110000101101) && ({row_reg, col_reg}<22'b0111010100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010100000001010111) && ({row_reg, col_reg}<22'b0111010100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010100000010000010) && ({row_reg, col_reg}<22'b0111010100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010100000111010111) && ({row_reg, col_reg}<22'b0111010100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111010100001000000010) && ({row_reg, col_reg}<22'b0111010100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010100001010000010) && ({row_reg, col_reg}<22'b0111010100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010100001010101101) && ({row_reg, col_reg}<22'b0111010100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010100010000000010) && ({row_reg, col_reg}<22'b0111010100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010100010000101101) && ({row_reg, col_reg}<22'b0111010100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010100100001010111) && ({row_reg, col_reg}<22'b0111010100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010100100010000010) && ({row_reg, col_reg}<22'b0111010100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010100100111010111) && ({row_reg, col_reg}<22'b0111010100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010100101000000010) && ({row_reg, col_reg}<22'b0111010100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010100101010000010) && ({row_reg, col_reg}<22'b0111010100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010100101010101101) && ({row_reg, col_reg}<22'b0111010100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010100110000000010) && ({row_reg, col_reg}<22'b0111010100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010100110000101101) && ({row_reg, col_reg}<22'b0111010101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010101000001010111) && ({row_reg, col_reg}<22'b0111010101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111010101000010000010) && ({row_reg, col_reg}<22'b0111010101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010101000111010111) && ({row_reg, col_reg}<22'b0111010101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010101001000000010) && ({row_reg, col_reg}<22'b0111010101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010101001010000010) && ({row_reg, col_reg}<22'b0111010101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010101001010101101) && ({row_reg, col_reg}<22'b0111010101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010101010000000010) && ({row_reg, col_reg}<22'b0111010101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010101010000101101) && ({row_reg, col_reg}<22'b0111010101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010101100001010111) && ({row_reg, col_reg}<22'b0111010101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111010101100010000010) && ({row_reg, col_reg}<22'b0111010101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010101100111010111) && ({row_reg, col_reg}<22'b0111010101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010101101000000010) && ({row_reg, col_reg}<22'b0111010101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010101101010000010) && ({row_reg, col_reg}<22'b0111010101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010101101010101101) && ({row_reg, col_reg}<22'b0111010101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010101110000000010) && ({row_reg, col_reg}<22'b0111010101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010101110000101101) && ({row_reg, col_reg}<22'b0111010110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010110000001010111) && ({row_reg, col_reg}<22'b0111010110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111010110000010000010) && ({row_reg, col_reg}<22'b0111010110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010110000111010111) && ({row_reg, col_reg}<22'b0111010110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010110001000000010) && ({row_reg, col_reg}<22'b0111010110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010110001010000010) && ({row_reg, col_reg}<22'b0111010110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010110001010101101) && ({row_reg, col_reg}<22'b0111010110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010110010000000010) && ({row_reg, col_reg}<22'b0111010110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010110010000101101) && ({row_reg, col_reg}<22'b0111010110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010110100001010111) && ({row_reg, col_reg}<22'b0111010110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010110100010000010) && ({row_reg, col_reg}<22'b0111010110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010110100111010111) && ({row_reg, col_reg}<22'b0111010110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010110101000000010) && ({row_reg, col_reg}<22'b0111010110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010110101010000010) && ({row_reg, col_reg}<22'b0111010110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010110101010101101) && ({row_reg, col_reg}<22'b0111010110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010110110000000010) && ({row_reg, col_reg}<22'b0111010110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010110110000101101) && ({row_reg, col_reg}<22'b0111010111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010111000001010111) && ({row_reg, col_reg}<22'b0111010111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111010111000010000010) && ({row_reg, col_reg}<22'b0111010111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010111000111010111) && ({row_reg, col_reg}<22'b0111010111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010111001000000010) && ({row_reg, col_reg}<22'b0111010111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010111001010000010) && ({row_reg, col_reg}<22'b0111010111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010111001010101101) && ({row_reg, col_reg}<22'b0111010111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010111010000000010) && ({row_reg, col_reg}<22'b0111010111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010111010000101101) && ({row_reg, col_reg}<22'b0111010111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010111100001010111) && ({row_reg, col_reg}<22'b0111010111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010111100010000010) && ({row_reg, col_reg}<22'b0111010111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111010111100111010111) && ({row_reg, col_reg}<22'b0111010111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111010111101000000010) && ({row_reg, col_reg}<22'b0111010111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010111101010000010) && ({row_reg, col_reg}<22'b0111010111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010111101010101101) && ({row_reg, col_reg}<22'b0111010111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111010111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111010111110000000010) && ({row_reg, col_reg}<22'b0111010111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111010111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111010111110000101101) && ({row_reg, col_reg}<22'b0111011000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011000000001010111) && ({row_reg, col_reg}<22'b0111011000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011000000010000010) && ({row_reg, col_reg}<22'b0111011000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011000000111010111) && ({row_reg, col_reg}<22'b0111011000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011000001000000010) && ({row_reg, col_reg}<22'b0111011000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011000001010000010) && ({row_reg, col_reg}<22'b0111011000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011000001010101101) && ({row_reg, col_reg}<22'b0111011000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011000010000000010) && ({row_reg, col_reg}<22'b0111011000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011000010000101101) && ({row_reg, col_reg}<22'b0111011000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011000100001010111) && ({row_reg, col_reg}<22'b0111011000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011000100010000010) && ({row_reg, col_reg}<22'b0111011000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011000100111010111) && ({row_reg, col_reg}<22'b0111011000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011000101000000010) && ({row_reg, col_reg}<22'b0111011000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011000101010000010) && ({row_reg, col_reg}<22'b0111011000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011000101010101101) && ({row_reg, col_reg}<22'b0111011000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011000110000000010) && ({row_reg, col_reg}<22'b0111011000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011000110000101101) && ({row_reg, col_reg}<22'b0111011001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011001000001010111) && ({row_reg, col_reg}<22'b0111011001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011001000010000010) && ({row_reg, col_reg}<22'b0111011001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011001000111010111) && ({row_reg, col_reg}<22'b0111011001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011001001000000010) && ({row_reg, col_reg}<22'b0111011001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011001001010000010) && ({row_reg, col_reg}<22'b0111011001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011001001010101101) && ({row_reg, col_reg}<22'b0111011001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011001010000000010) && ({row_reg, col_reg}<22'b0111011001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011001010000101101) && ({row_reg, col_reg}<22'b0111011001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011001100001010111) && ({row_reg, col_reg}<22'b0111011001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011001100010000010) && ({row_reg, col_reg}<22'b0111011001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011001100111010111) && ({row_reg, col_reg}<22'b0111011001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011001101000000010) && ({row_reg, col_reg}<22'b0111011001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011001101010000010) && ({row_reg, col_reg}<22'b0111011001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011001101010101101) && ({row_reg, col_reg}<22'b0111011001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011001110000000010) && ({row_reg, col_reg}<22'b0111011001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011001110000101101) && ({row_reg, col_reg}<22'b0111011010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011010000001010111) && ({row_reg, col_reg}<22'b0111011010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011010000010000010) && ({row_reg, col_reg}<22'b0111011010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011010000111010111) && ({row_reg, col_reg}<22'b0111011010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011010001000000010) && ({row_reg, col_reg}<22'b0111011010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011010001010000010) && ({row_reg, col_reg}<22'b0111011010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011010001010101101) && ({row_reg, col_reg}<22'b0111011010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011010010000000010) && ({row_reg, col_reg}<22'b0111011010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011010010000101101) && ({row_reg, col_reg}<22'b0111011010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011010100001010111) && ({row_reg, col_reg}<22'b0111011010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011010100010000010) && ({row_reg, col_reg}<22'b0111011010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011010100111010111) && ({row_reg, col_reg}<22'b0111011010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011010101000000010) && ({row_reg, col_reg}<22'b0111011010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011010101010000010) && ({row_reg, col_reg}<22'b0111011010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011010101010101101) && ({row_reg, col_reg}<22'b0111011010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011010110000000010) && ({row_reg, col_reg}<22'b0111011010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011010110000101101) && ({row_reg, col_reg}<22'b0111011011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011011000001010111) && ({row_reg, col_reg}<22'b0111011011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011011000010000010) && ({row_reg, col_reg}<22'b0111011011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011011000111010111) && ({row_reg, col_reg}<22'b0111011011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011011001000000010) && ({row_reg, col_reg}<22'b0111011011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011011001010000010) && ({row_reg, col_reg}<22'b0111011011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011011001010101101) && ({row_reg, col_reg}<22'b0111011011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011011010000000010) && ({row_reg, col_reg}<22'b0111011011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011011010000101101) && ({row_reg, col_reg}<22'b0111011011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011011100001010111) && ({row_reg, col_reg}<22'b0111011011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011011100010000010) && ({row_reg, col_reg}<22'b0111011011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011011100111010111) && ({row_reg, col_reg}<22'b0111011011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011011101000000010) && ({row_reg, col_reg}<22'b0111011011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011011101010000010) && ({row_reg, col_reg}<22'b0111011011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011011101010101101) && ({row_reg, col_reg}<22'b0111011011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011011110000000010) && ({row_reg, col_reg}<22'b0111011011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011011110000101101) && ({row_reg, col_reg}<22'b0111011100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011100000001010111) && ({row_reg, col_reg}<22'b0111011100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011100000010000010) && ({row_reg, col_reg}<22'b0111011100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011100000111010111) && ({row_reg, col_reg}<22'b0111011100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111011100001000000010) && ({row_reg, col_reg}<22'b0111011100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011100001010000010) && ({row_reg, col_reg}<22'b0111011100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011100001010101101) && ({row_reg, col_reg}<22'b0111011100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011100010000000010) && ({row_reg, col_reg}<22'b0111011100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011100010000101101) && ({row_reg, col_reg}<22'b0111011100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011100100001010111) && ({row_reg, col_reg}<22'b0111011100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011100100010000010) && ({row_reg, col_reg}<22'b0111011100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011100100111010111) && ({row_reg, col_reg}<22'b0111011100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111011100101000000010) && ({row_reg, col_reg}<22'b0111011100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011100101010000010) && ({row_reg, col_reg}<22'b0111011100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011100101010101101) && ({row_reg, col_reg}<22'b0111011100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011100110000000010) && ({row_reg, col_reg}<22'b0111011100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011100110000101101) && ({row_reg, col_reg}<22'b0111011101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011101000001010111) && ({row_reg, col_reg}<22'b0111011101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011101000010000010) && ({row_reg, col_reg}<22'b0111011101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011101000111010111) && ({row_reg, col_reg}<22'b0111011101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111011101001000000010) && ({row_reg, col_reg}<22'b0111011101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011101001010000010) && ({row_reg, col_reg}<22'b0111011101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011101001010101101) && ({row_reg, col_reg}<22'b0111011101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011101010000000010) && ({row_reg, col_reg}<22'b0111011101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011101010000101101) && ({row_reg, col_reg}<22'b0111011101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011101100001010111) && ({row_reg, col_reg}<22'b0111011101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011101100010000010) && ({row_reg, col_reg}<22'b0111011101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011101100111010111) && ({row_reg, col_reg}<22'b0111011101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111011101101000000010) && ({row_reg, col_reg}<22'b0111011101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011101101010000010) && ({row_reg, col_reg}<22'b0111011101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011101101010101101) && ({row_reg, col_reg}<22'b0111011101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011101110000000010) && ({row_reg, col_reg}<22'b0111011101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011101110000101101) && ({row_reg, col_reg}<22'b0111011110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011110000001010111) && ({row_reg, col_reg}<22'b0111011110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111011110000010000010) && ({row_reg, col_reg}<22'b0111011110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011110000111010111) && ({row_reg, col_reg}<22'b0111011110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111011110001000000010) && ({row_reg, col_reg}<22'b0111011110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011110001010000010) && ({row_reg, col_reg}<22'b0111011110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011110001010101101) && ({row_reg, col_reg}<22'b0111011110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011110010000000010) && ({row_reg, col_reg}<22'b0111011110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011110010000101101) && ({row_reg, col_reg}<22'b0111011110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011110100001010111) && ({row_reg, col_reg}<22'b0111011110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111011110100010000010) && ({row_reg, col_reg}<22'b0111011110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011110100111010111) && ({row_reg, col_reg}<22'b0111011110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111011110101000000010) && ({row_reg, col_reg}<22'b0111011110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011110101010000010) && ({row_reg, col_reg}<22'b0111011110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011110101010101101) && ({row_reg, col_reg}<22'b0111011110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011110110000000010) && ({row_reg, col_reg}<22'b0111011110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011110110000101101) && ({row_reg, col_reg}<22'b0111011111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011111000001010111) && ({row_reg, col_reg}<22'b0111011111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111011111000010000010) && ({row_reg, col_reg}<22'b0111011111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011111000111010111) && ({row_reg, col_reg}<22'b0111011111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111011111001000000010) && ({row_reg, col_reg}<22'b0111011111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011111001010000010) && ({row_reg, col_reg}<22'b0111011111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011111001010101101) && ({row_reg, col_reg}<22'b0111011111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011111010000000010) && ({row_reg, col_reg}<22'b0111011111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011111010000101101) && ({row_reg, col_reg}<22'b0111011111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011111100001010111) && ({row_reg, col_reg}<22'b0111011111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111011111100010000010) && ({row_reg, col_reg}<22'b0111011111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111011111100111010111) && ({row_reg, col_reg}<22'b0111011111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111011111101000000010) && ({row_reg, col_reg}<22'b0111011111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011111101010000010) && ({row_reg, col_reg}<22'b0111011111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011111101010101101) && ({row_reg, col_reg}<22'b0111011111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111011111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111011111110000000010) && ({row_reg, col_reg}<22'b0111011111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111011111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111011111110000101101) && ({row_reg, col_reg}<22'b0111100000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100000000001010111) && ({row_reg, col_reg}<22'b0111100000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111100000000010000010) && ({row_reg, col_reg}<22'b0111100000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100000000111010111) && ({row_reg, col_reg}<22'b0111100000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100000001000000010) && ({row_reg, col_reg}<22'b0111100000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100000001010000010) && ({row_reg, col_reg}<22'b0111100000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100000001010101101) && ({row_reg, col_reg}<22'b0111100000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100000010000000010) && ({row_reg, col_reg}<22'b0111100000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100000010000101101) && ({row_reg, col_reg}<22'b0111100000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100000100001010111) && ({row_reg, col_reg}<22'b0111100000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111100000100010000010) && ({row_reg, col_reg}<22'b0111100000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100000100111010111) && ({row_reg, col_reg}<22'b0111100000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100000101000000010) && ({row_reg, col_reg}<22'b0111100000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100000101010000010) && ({row_reg, col_reg}<22'b0111100000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100000101010101101) && ({row_reg, col_reg}<22'b0111100000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100000110000000010) && ({row_reg, col_reg}<22'b0111100000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100000110000101101) && ({row_reg, col_reg}<22'b0111100001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100001000001010111) && ({row_reg, col_reg}<22'b0111100001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111100001000010000010) && ({row_reg, col_reg}<22'b0111100001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100001000111010111) && ({row_reg, col_reg}<22'b0111100001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100001001000000010) && ({row_reg, col_reg}<22'b0111100001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100001001010000010) && ({row_reg, col_reg}<22'b0111100001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100001001010101101) && ({row_reg, col_reg}<22'b0111100001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100001010000000010) && ({row_reg, col_reg}<22'b0111100001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100001010000101101) && ({row_reg, col_reg}<22'b0111100001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100001100001010111) && ({row_reg, col_reg}<22'b0111100001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100001100010000010) && ({row_reg, col_reg}<22'b0111100001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100001100111010111) && ({row_reg, col_reg}<22'b0111100001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100001101000000010) && ({row_reg, col_reg}<22'b0111100001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100001101010000010) && ({row_reg, col_reg}<22'b0111100001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100001101010101101) && ({row_reg, col_reg}<22'b0111100001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100001110000000010) && ({row_reg, col_reg}<22'b0111100001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100001110000101101) && ({row_reg, col_reg}<22'b0111100010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100010000001010111) && ({row_reg, col_reg}<22'b0111100010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100010000010000010) && ({row_reg, col_reg}<22'b0111100010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100010000111010111) && ({row_reg, col_reg}<22'b0111100010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100010001000000010) && ({row_reg, col_reg}<22'b0111100010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100010001010000010) && ({row_reg, col_reg}<22'b0111100010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100010001010101101) && ({row_reg, col_reg}<22'b0111100010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100010010000000010) && ({row_reg, col_reg}<22'b0111100010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100010010000101101) && ({row_reg, col_reg}<22'b0111100010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100010100001010111) && ({row_reg, col_reg}<22'b0111100010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100010100010000010) && ({row_reg, col_reg}<22'b0111100010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100010100111010111) && ({row_reg, col_reg}<22'b0111100010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100010101000000010) && ({row_reg, col_reg}<22'b0111100010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100010101010000010) && ({row_reg, col_reg}<22'b0111100010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100010101010101101) && ({row_reg, col_reg}<22'b0111100010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100010110000000010) && ({row_reg, col_reg}<22'b0111100010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100010110000101101) && ({row_reg, col_reg}<22'b0111100011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100011000001010111) && ({row_reg, col_reg}<22'b0111100011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100011000010000010) && ({row_reg, col_reg}<22'b0111100011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100011000111010111) && ({row_reg, col_reg}<22'b0111100011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100011001000000010) && ({row_reg, col_reg}<22'b0111100011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100011001010000010) && ({row_reg, col_reg}<22'b0111100011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100011001010101101) && ({row_reg, col_reg}<22'b0111100011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100011010000000010) && ({row_reg, col_reg}<22'b0111100011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100011010000101101) && ({row_reg, col_reg}<22'b0111100011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100011100001010111) && ({row_reg, col_reg}<22'b0111100011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100011100010000010) && ({row_reg, col_reg}<22'b0111100011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100011100111010111) && ({row_reg, col_reg}<22'b0111100011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100011101000000010) && ({row_reg, col_reg}<22'b0111100011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100011101010000010) && ({row_reg, col_reg}<22'b0111100011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100011101010101101) && ({row_reg, col_reg}<22'b0111100011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100011110000000010) && ({row_reg, col_reg}<22'b0111100011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100011110000101101) && ({row_reg, col_reg}<22'b0111100100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100100000001010111) && ({row_reg, col_reg}<22'b0111100100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100100000010000010) && ({row_reg, col_reg}<22'b0111100100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100100000111010111) && ({row_reg, col_reg}<22'b0111100100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100100001000000010) && ({row_reg, col_reg}<22'b0111100100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100100001010000010) && ({row_reg, col_reg}<22'b0111100100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100100001010101101) && ({row_reg, col_reg}<22'b0111100100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100100010000000010) && ({row_reg, col_reg}<22'b0111100100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100100010000101101) && ({row_reg, col_reg}<22'b0111100100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100100100001010111) && ({row_reg, col_reg}<22'b0111100100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100100100010000010) && ({row_reg, col_reg}<22'b0111100100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100100100111010111) && ({row_reg, col_reg}<22'b0111100100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100100101000000010) && ({row_reg, col_reg}<22'b0111100100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100100101010000010) && ({row_reg, col_reg}<22'b0111100100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100100101010101101) && ({row_reg, col_reg}<22'b0111100100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100100110000000010) && ({row_reg, col_reg}<22'b0111100100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100100110000101101) && ({row_reg, col_reg}<22'b0111100101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100101000001010111) && ({row_reg, col_reg}<22'b0111100101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100101000010000010) && ({row_reg, col_reg}<22'b0111100101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100101000111010111) && ({row_reg, col_reg}<22'b0111100101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100101001000000010) && ({row_reg, col_reg}<22'b0111100101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100101001010000010) && ({row_reg, col_reg}<22'b0111100101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100101001010101101) && ({row_reg, col_reg}<22'b0111100101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100101010000000010) && ({row_reg, col_reg}<22'b0111100101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100101010000101101) && ({row_reg, col_reg}<22'b0111100101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100101100001010111) && ({row_reg, col_reg}<22'b0111100101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100101100010000010) && ({row_reg, col_reg}<22'b0111100101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100101100111010111) && ({row_reg, col_reg}<22'b0111100101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100101101000000010) && ({row_reg, col_reg}<22'b0111100101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100101101010000010) && ({row_reg, col_reg}<22'b0111100101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100101101010101101) && ({row_reg, col_reg}<22'b0111100101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100101110000000010) && ({row_reg, col_reg}<22'b0111100101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100101110000101101) && ({row_reg, col_reg}<22'b0111100110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100110000001010111) && ({row_reg, col_reg}<22'b0111100110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100110000010000010) && ({row_reg, col_reg}<22'b0111100110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100110000111010111) && ({row_reg, col_reg}<22'b0111100110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111100110001000000010) && ({row_reg, col_reg}<22'b0111100110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100110001010000010) && ({row_reg, col_reg}<22'b0111100110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100110001010101101) && ({row_reg, col_reg}<22'b0111100110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100110010000000010) && ({row_reg, col_reg}<22'b0111100110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100110010000101101) && ({row_reg, col_reg}<22'b0111100110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100110100001010111) && ({row_reg, col_reg}<22'b0111100110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100110100010000010) && ({row_reg, col_reg}<22'b0111100110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100110100111010111) && ({row_reg, col_reg}<22'b0111100110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111100110101000000010) && ({row_reg, col_reg}<22'b0111100110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100110101010000010) && ({row_reg, col_reg}<22'b0111100110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100110101010101101) && ({row_reg, col_reg}<22'b0111100110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100110110000000010) && ({row_reg, col_reg}<22'b0111100110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100110110000101101) && ({row_reg, col_reg}<22'b0111100111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100111000001010111) && ({row_reg, col_reg}<22'b0111100111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100111000010000010) && ({row_reg, col_reg}<22'b0111100111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100111000111010111) && ({row_reg, col_reg}<22'b0111100111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111100111001000000010) && ({row_reg, col_reg}<22'b0111100111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100111001010000010) && ({row_reg, col_reg}<22'b0111100111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100111001010101101) && ({row_reg, col_reg}<22'b0111100111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100111010000000010) && ({row_reg, col_reg}<22'b0111100111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100111010000101101) && ({row_reg, col_reg}<22'b0111100111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100111100001010111) && ({row_reg, col_reg}<22'b0111100111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111100111100010000010) && ({row_reg, col_reg}<22'b0111100111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111100111100111010111) && ({row_reg, col_reg}<22'b0111100111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111100111101000000010) && ({row_reg, col_reg}<22'b0111100111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100111101010000010) && ({row_reg, col_reg}<22'b0111100111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100111101010101101) && ({row_reg, col_reg}<22'b0111100111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111100111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111100111110000000010) && ({row_reg, col_reg}<22'b0111100111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111100111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111100111110000101101) && ({row_reg, col_reg}<22'b0111101000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101000000001010111) && ({row_reg, col_reg}<22'b0111101000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111101000000010000010) && ({row_reg, col_reg}<22'b0111101000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101000000111010111) && ({row_reg, col_reg}<22'b0111101000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111101000001000000010) && ({row_reg, col_reg}<22'b0111101000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101000001010000010) && ({row_reg, col_reg}<22'b0111101000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101000001010101101) && ({row_reg, col_reg}<22'b0111101000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101000010000000010) && ({row_reg, col_reg}<22'b0111101000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101000010000101101) && ({row_reg, col_reg}<22'b0111101000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101000100001010111) && ({row_reg, col_reg}<22'b0111101000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111101000100010000010) && ({row_reg, col_reg}<22'b0111101000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101000100111010111) && ({row_reg, col_reg}<22'b0111101000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111101000101000000010) && ({row_reg, col_reg}<22'b0111101000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101000101010000010) && ({row_reg, col_reg}<22'b0111101000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101000101010101101) && ({row_reg, col_reg}<22'b0111101000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101000110000000010) && ({row_reg, col_reg}<22'b0111101000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101000110000101101) && ({row_reg, col_reg}<22'b0111101001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101001000001010111) && ({row_reg, col_reg}<22'b0111101001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111101001000010000010) && ({row_reg, col_reg}<22'b0111101001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101001000111010111) && ({row_reg, col_reg}<22'b0111101001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111101001001000000010) && ({row_reg, col_reg}<22'b0111101001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101001001010000010) && ({row_reg, col_reg}<22'b0111101001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101001001010101101) && ({row_reg, col_reg}<22'b0111101001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101001010000000010) && ({row_reg, col_reg}<22'b0111101001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101001010000101101) && ({row_reg, col_reg}<22'b0111101001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101001100001010111) && ({row_reg, col_reg}<22'b0111101001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111101001100010000010) && ({row_reg, col_reg}<22'b0111101001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101001100111010111) && ({row_reg, col_reg}<22'b0111101001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101001101000000010) && ({row_reg, col_reg}<22'b0111101001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101001101010000010) && ({row_reg, col_reg}<22'b0111101001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101001101010101101) && ({row_reg, col_reg}<22'b0111101001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101001110000000010) && ({row_reg, col_reg}<22'b0111101001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101001110000101101) && ({row_reg, col_reg}<22'b0111101010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101010000001010111) && ({row_reg, col_reg}<22'b0111101010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111101010000010000010) && ({row_reg, col_reg}<22'b0111101010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101010000111010111) && ({row_reg, col_reg}<22'b0111101010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101010001000000010) && ({row_reg, col_reg}<22'b0111101010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101010001010000010) && ({row_reg, col_reg}<22'b0111101010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101010001010101101) && ({row_reg, col_reg}<22'b0111101010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101010010000000010) && ({row_reg, col_reg}<22'b0111101010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101010010000101101) && ({row_reg, col_reg}<22'b0111101010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101010100001010111) && ({row_reg, col_reg}<22'b0111101010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111101010100010000010) && ({row_reg, col_reg}<22'b0111101010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101010100111010111) && ({row_reg, col_reg}<22'b0111101010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101010101000000010) && ({row_reg, col_reg}<22'b0111101010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101010101010000010) && ({row_reg, col_reg}<22'b0111101010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101010101010101101) && ({row_reg, col_reg}<22'b0111101010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101010110000000010) && ({row_reg, col_reg}<22'b0111101010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101010110000101101) && ({row_reg, col_reg}<22'b0111101011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101011000001010111) && ({row_reg, col_reg}<22'b0111101011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111101011000010000010) && ({row_reg, col_reg}<22'b0111101011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101011000111010111) && ({row_reg, col_reg}<22'b0111101011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101011001000000010) && ({row_reg, col_reg}<22'b0111101011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101011001010000010) && ({row_reg, col_reg}<22'b0111101011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101011001010101101) && ({row_reg, col_reg}<22'b0111101011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101011010000000010) && ({row_reg, col_reg}<22'b0111101011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101011010000101101) && ({row_reg, col_reg}<22'b0111101011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101011100001010111) && ({row_reg, col_reg}<22'b0111101011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101011100010000010) && ({row_reg, col_reg}<22'b0111101011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101011100111010111) && ({row_reg, col_reg}<22'b0111101011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101011101000000010) && ({row_reg, col_reg}<22'b0111101011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101011101010000010) && ({row_reg, col_reg}<22'b0111101011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101011101010101101) && ({row_reg, col_reg}<22'b0111101011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101011110000000010) && ({row_reg, col_reg}<22'b0111101011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101011110000101101) && ({row_reg, col_reg}<22'b0111101100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101100000001010111) && ({row_reg, col_reg}<22'b0111101100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101100000010000010) && ({row_reg, col_reg}<22'b0111101100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101100000111010111) && ({row_reg, col_reg}<22'b0111101100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101100001000000010) && ({row_reg, col_reg}<22'b0111101100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101100001010000010) && ({row_reg, col_reg}<22'b0111101100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101100001010101101) && ({row_reg, col_reg}<22'b0111101100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101100010000000010) && ({row_reg, col_reg}<22'b0111101100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101100010000101101) && ({row_reg, col_reg}<22'b0111101100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101100100001010111) && ({row_reg, col_reg}<22'b0111101100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101100100010000010) && ({row_reg, col_reg}<22'b0111101100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101100100111010111) && ({row_reg, col_reg}<22'b0111101100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101100101000000010) && ({row_reg, col_reg}<22'b0111101100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101100101010000010) && ({row_reg, col_reg}<22'b0111101100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101100101010101101) && ({row_reg, col_reg}<22'b0111101100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101100110000000010) && ({row_reg, col_reg}<22'b0111101100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101100110000101101) && ({row_reg, col_reg}<22'b0111101101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101101000001010111) && ({row_reg, col_reg}<22'b0111101101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101101000010000010) && ({row_reg, col_reg}<22'b0111101101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101101000111010111) && ({row_reg, col_reg}<22'b0111101101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101101001000000010) && ({row_reg, col_reg}<22'b0111101101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101101001010000010) && ({row_reg, col_reg}<22'b0111101101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101101001010101101) && ({row_reg, col_reg}<22'b0111101101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101101010000000010) && ({row_reg, col_reg}<22'b0111101101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101101010000101101) && ({row_reg, col_reg}<22'b0111101101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101101100001010111) && ({row_reg, col_reg}<22'b0111101101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101101100010000010) && ({row_reg, col_reg}<22'b0111101101100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101101100111010111) && ({row_reg, col_reg}<22'b0111101101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101101101000000010) && ({row_reg, col_reg}<22'b0111101101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101101101010000010) && ({row_reg, col_reg}<22'b0111101101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101101101010101101) && ({row_reg, col_reg}<22'b0111101101110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101101110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101101110000000010) && ({row_reg, col_reg}<22'b0111101101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101101110000101101) && ({row_reg, col_reg}<22'b0111101110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101110000001010111) && ({row_reg, col_reg}<22'b0111101110000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101110000010000010) && ({row_reg, col_reg}<22'b0111101110000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101110000111010111) && ({row_reg, col_reg}<22'b0111101110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101110001000000010) && ({row_reg, col_reg}<22'b0111101110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101110001010000010) && ({row_reg, col_reg}<22'b0111101110001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101110001010101101) && ({row_reg, col_reg}<22'b0111101110010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101110010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101110010000000010) && ({row_reg, col_reg}<22'b0111101110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101110010000101101) && ({row_reg, col_reg}<22'b0111101110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101110100001010111) && ({row_reg, col_reg}<22'b0111101110100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101110100010000010) && ({row_reg, col_reg}<22'b0111101110100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101110100111010111) && ({row_reg, col_reg}<22'b0111101110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101110101000000010) && ({row_reg, col_reg}<22'b0111101110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101110101010000010) && ({row_reg, col_reg}<22'b0111101110101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101110101010101101) && ({row_reg, col_reg}<22'b0111101110110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101110110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101110110000000010) && ({row_reg, col_reg}<22'b0111101110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101110110000101101) && ({row_reg, col_reg}<22'b0111101111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101111000001010111) && ({row_reg, col_reg}<22'b0111101111000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101111000010000010) && ({row_reg, col_reg}<22'b0111101111000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101111000111010111) && ({row_reg, col_reg}<22'b0111101111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101111001000000010) && ({row_reg, col_reg}<22'b0111101111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101111001010000010) && ({row_reg, col_reg}<22'b0111101111001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101111001010101101) && ({row_reg, col_reg}<22'b0111101111010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101111010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101111010000000010) && ({row_reg, col_reg}<22'b0111101111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101111010000101101) && ({row_reg, col_reg}<22'b0111101111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101111100001010111) && ({row_reg, col_reg}<22'b0111101111100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101111100010000010) && ({row_reg, col_reg}<22'b0111101111100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111101111100111010111) && ({row_reg, col_reg}<22'b0111101111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111101111101000000010) && ({row_reg, col_reg}<22'b0111101111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101111101010000010) && ({row_reg, col_reg}<22'b0111101111101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101111101010101101) && ({row_reg, col_reg}<22'b0111101111110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111101111110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111101111110000000010) && ({row_reg, col_reg}<22'b0111101111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111101111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111101111110000101101) && ({row_reg, col_reg}<22'b0111110000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110000000001010111) && ({row_reg, col_reg}<22'b0111110000000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110000000010000010) && ({row_reg, col_reg}<22'b0111110000000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110000000111010111) && ({row_reg, col_reg}<22'b0111110000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110000001000000010) && ({row_reg, col_reg}<22'b0111110000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110000001010000010) && ({row_reg, col_reg}<22'b0111110000001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110000001010101101) && ({row_reg, col_reg}<22'b0111110000010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110000010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110000010000000010) && ({row_reg, col_reg}<22'b0111110000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110000010000101101) && ({row_reg, col_reg}<22'b0111110000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110000100001010111) && ({row_reg, col_reg}<22'b0111110000100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110000100010000010) && ({row_reg, col_reg}<22'b0111110000100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110000100111010111) && ({row_reg, col_reg}<22'b0111110000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110000101000000010) && ({row_reg, col_reg}<22'b0111110000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110000101010000010) && ({row_reg, col_reg}<22'b0111110000101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110000101010101101) && ({row_reg, col_reg}<22'b0111110000110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110000110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110000110000000010) && ({row_reg, col_reg}<22'b0111110000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110000110000101101) && ({row_reg, col_reg}<22'b0111110001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110001000001010111) && ({row_reg, col_reg}<22'b0111110001000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001000010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110001000010000010) && ({row_reg, col_reg}<22'b0111110001000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110001000111010111) && ({row_reg, col_reg}<22'b0111110001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110001001000000010) && ({row_reg, col_reg}<22'b0111110001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110001001010000010) && ({row_reg, col_reg}<22'b0111110001001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110001001010101101) && ({row_reg, col_reg}<22'b0111110001010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110001010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110001010000000010) && ({row_reg, col_reg}<22'b0111110001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110001010000101101) && ({row_reg, col_reg}<22'b0111110001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110001100001010111) && ({row_reg, col_reg}<22'b0111110001100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001100010000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110001100010000010) && ({row_reg, col_reg}<22'b0111110001100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110001100111010111) && ({row_reg, col_reg}<22'b0111110001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110001101000000010) && ({row_reg, col_reg}<22'b0111110001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110001101010000010) && ({row_reg, col_reg}<22'b0111110001101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110001101010101101) && ({row_reg, col_reg}<22'b0111110001110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110001110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110001110000000010) && ({row_reg, col_reg}<22'b0111110001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110001110000101101) && ({row_reg, col_reg}<22'b0111110010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110010000001010111) && ({row_reg, col_reg}<22'b0111110010000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110010000010000010) && ({row_reg, col_reg}<22'b0111110010000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110010000111010111) && ({row_reg, col_reg}<22'b0111110010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110010001000000010) && ({row_reg, col_reg}<22'b0111110010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110010001010000010) && ({row_reg, col_reg}<22'b0111110010001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110010001010101101) && ({row_reg, col_reg}<22'b0111110010010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110010010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110010010000000010) && ({row_reg, col_reg}<22'b0111110010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110010010000101101) && ({row_reg, col_reg}<22'b0111110010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110010100001010111) && ({row_reg, col_reg}<22'b0111110010100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110010100010000010) && ({row_reg, col_reg}<22'b0111110010100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110010100111010111) && ({row_reg, col_reg}<22'b0111110010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110010101000000010) && ({row_reg, col_reg}<22'b0111110010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110010101010000010) && ({row_reg, col_reg}<22'b0111110010101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110010101010101101) && ({row_reg, col_reg}<22'b0111110010110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110010110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110010110000000010) && ({row_reg, col_reg}<22'b0111110010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110010110000101101) && ({row_reg, col_reg}<22'b0111110011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110011000001010111) && ({row_reg, col_reg}<22'b0111110011000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110011000010000010) && ({row_reg, col_reg}<22'b0111110011000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110011000111010111) && ({row_reg, col_reg}<22'b0111110011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110011001000000010) && ({row_reg, col_reg}<22'b0111110011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110011001010000010) && ({row_reg, col_reg}<22'b0111110011001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110011001010101101) && ({row_reg, col_reg}<22'b0111110011010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110011010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110011010000000010) && ({row_reg, col_reg}<22'b0111110011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110011010000101101) && ({row_reg, col_reg}<22'b0111110011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110011100001010111) && ({row_reg, col_reg}<22'b0111110011100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011100010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110011100010000010) && ({row_reg, col_reg}<22'b0111110011100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110011100111010111) && ({row_reg, col_reg}<22'b0111110011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110011101000000010) && ({row_reg, col_reg}<22'b0111110011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110011101010000010) && ({row_reg, col_reg}<22'b0111110011101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110011101010101101) && ({row_reg, col_reg}<22'b0111110011110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110011110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110011110000000010) && ({row_reg, col_reg}<22'b0111110011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110011110000101101) && ({row_reg, col_reg}<22'b0111110100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110100000001010111) && ({row_reg, col_reg}<22'b0111110100000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100000010000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110100000010000010) && ({row_reg, col_reg}<22'b0111110100000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110100000111010111) && ({row_reg, col_reg}<22'b0111110100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110100001000000010) && ({row_reg, col_reg}<22'b0111110100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110100001010000010) && ({row_reg, col_reg}<22'b0111110100001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110100001010101101) && ({row_reg, col_reg}<22'b0111110100010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110100010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110100010000000010) && ({row_reg, col_reg}<22'b0111110100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110100010000101101) && ({row_reg, col_reg}<22'b0111110100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110100100001010111) && ({row_reg, col_reg}<22'b0111110100100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100100010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110100100010000010) && ({row_reg, col_reg}<22'b0111110100100111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110100100111010111) && ({row_reg, col_reg}<22'b0111110100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110100101000000010) && ({row_reg, col_reg}<22'b0111110100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110100101010000010) && ({row_reg, col_reg}<22'b0111110100101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100101010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110100101010101101) && ({row_reg, col_reg}<22'b0111110100110000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110100110000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110100110000000010) && ({row_reg, col_reg}<22'b0111110100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110100110000101101) && ({row_reg, col_reg}<22'b0111110101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110101000001010111) && ({row_reg, col_reg}<22'b0111110101000010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101000010000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111110101000010000010) && ({row_reg, col_reg}<22'b0111110101000111010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110101000111010111) && ({row_reg, col_reg}<22'b0111110101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101001000000010) && ({row_reg, col_reg}<22'b0111110101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110101001010000010) && ({row_reg, col_reg}<22'b0111110101001010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101001010101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110101001010101101) && ({row_reg, col_reg}<22'b0111110101010000000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110101010000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110101010000000010) && ({row_reg, col_reg}<22'b0111110101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110101010000101101) && ({row_reg, col_reg}<22'b0111110101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110101100001010111) && ({row_reg, col_reg}<22'b0111110101100010000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101100010000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b0111110101100010000010) && ({row_reg, col_reg}<22'b0111110101100010001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100010001110) && ({row_reg, col_reg}<22'b0111110101100010010101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100010010101) && ({row_reg, col_reg}<22'b0111110101100010100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100010100010) && ({row_reg, col_reg}<22'b0111110101100010101001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100010101001) && ({row_reg, col_reg}<22'b0111110101100010110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100010110110) && ({row_reg, col_reg}<22'b0111110101100010111101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100010111101) && ({row_reg, col_reg}<22'b0111110101100011001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100011001010) && ({row_reg, col_reg}<22'b0111110101100011010001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100011010001) && ({row_reg, col_reg}<22'b0111110101100011011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100011011110) && ({row_reg, col_reg}<22'b0111110101100011100101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100011100101) && ({row_reg, col_reg}<22'b0111110101100011110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100011110010) && ({row_reg, col_reg}<22'b0111110101100011111001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100011111001) && ({row_reg, col_reg}<22'b0111110101100100000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100100000110) && ({row_reg, col_reg}<22'b0111110101100100001101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100100001101) && ({row_reg, col_reg}<22'b0111110101100100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100100011010) && ({row_reg, col_reg}<22'b0111110101100100100001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100100100001) && ({row_reg, col_reg}<22'b0111110101100100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100100101110) && ({row_reg, col_reg}<22'b0111110101100100110101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100100110101) && ({row_reg, col_reg}<22'b0111110101100101000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100101000010) && ({row_reg, col_reg}<22'b0111110101100101001001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100101001001) && ({row_reg, col_reg}<22'b0111110101100101010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100101010110) && ({row_reg, col_reg}<22'b0111110101100101011101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100101011101) && ({row_reg, col_reg}<22'b0111110101100101101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100101101010) && ({row_reg, col_reg}<22'b0111110101100101110001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100101110001) && ({row_reg, col_reg}<22'b0111110101100101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100101111110) && ({row_reg, col_reg}<22'b0111110101100110000101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100110000101) && ({row_reg, col_reg}<22'b0111110101100110010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100110010010) && ({row_reg, col_reg}<22'b0111110101100110011001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100110011001) && ({row_reg, col_reg}<22'b0111110101100110100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100110100110) && ({row_reg, col_reg}<22'b0111110101100110101101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100110101101) && ({row_reg, col_reg}<22'b0111110101100110111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100110111010) && ({row_reg, col_reg}<22'b0111110101100111000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100111000001) && ({row_reg, col_reg}<22'b0111110101100111001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100111001110) && ({row_reg, col_reg}<22'b0111110101100111010101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101100111010101) && ({row_reg, col_reg}<22'b0111110101100111010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101100111010111) && ({row_reg, col_reg}<22'b0111110101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101000000010) && ({row_reg, col_reg}<22'b0111110101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110101101010000010) && ({row_reg, col_reg}<22'b0111110101101010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101101010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0111110101101010101101) && ({row_reg, col_reg}<22'b0111110101101010110001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101010110001) && ({row_reg, col_reg}<22'b0111110101101010111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101010111110) && ({row_reg, col_reg}<22'b0111110101101011000101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101011000101) && ({row_reg, col_reg}<22'b0111110101101011010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101011010010) && ({row_reg, col_reg}<22'b0111110101101011011001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101011011001) && ({row_reg, col_reg}<22'b0111110101101011100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101011100110) && ({row_reg, col_reg}<22'b0111110101101011101101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101011101101) && ({row_reg, col_reg}<22'b0111110101101011111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101011111010) && ({row_reg, col_reg}<22'b0111110101101100000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101100000001) && ({row_reg, col_reg}<22'b0111110101101100001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101100001110) && ({row_reg, col_reg}<22'b0111110101101100010101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101100010101) && ({row_reg, col_reg}<22'b0111110101101100100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101100100010) && ({row_reg, col_reg}<22'b0111110101101100101001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101100101001) && ({row_reg, col_reg}<22'b0111110101101100110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101100110110) && ({row_reg, col_reg}<22'b0111110101101100111101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101100111101) && ({row_reg, col_reg}<22'b0111110101101101001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101101001010) && ({row_reg, col_reg}<22'b0111110101101101010001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101101010001) && ({row_reg, col_reg}<22'b0111110101101101011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101101011110) && ({row_reg, col_reg}<22'b0111110101101101100101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101101100101) && ({row_reg, col_reg}<22'b0111110101101101110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101101110010) && ({row_reg, col_reg}<22'b0111110101101101111001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101101111001) && ({row_reg, col_reg}<22'b0111110101101110000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101110000110) && ({row_reg, col_reg}<22'b0111110101101110001101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101110001101) && ({row_reg, col_reg}<22'b0111110101101110011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101110011010) && ({row_reg, col_reg}<22'b0111110101101110100001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101110100001) && ({row_reg, col_reg}<22'b0111110101101110101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101110101110) && ({row_reg, col_reg}<22'b0111110101101110110101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101110110101) && ({row_reg, col_reg}<22'b0111110101101111000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101111000010) && ({row_reg, col_reg}<22'b0111110101101111001001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101111001001) && ({row_reg, col_reg}<22'b0111110101101111010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101111010110) && ({row_reg, col_reg}<22'b0111110101101111011101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101111011101) && ({row_reg, col_reg}<22'b0111110101101111101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101111101010) && ({row_reg, col_reg}<22'b0111110101101111110001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111110101101111110001) && ({row_reg, col_reg}<22'b0111110101101111111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110101101111111110) && ({row_reg, col_reg}<22'b0111110101110000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==22'b0111110101110000000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b0111110101110000000010) && ({row_reg, col_reg}<22'b0111110101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110101110000101101) && ({row_reg, col_reg}<22'b0111110110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110110000001010111) && ({row_reg, col_reg}<22'b0111110110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110110001000000010) && ({row_reg, col_reg}<22'b0111110110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110110001010000010) && ({row_reg, col_reg}<22'b0111110110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110110010000101101) && ({row_reg, col_reg}<22'b0111110110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110110100001010111) && ({row_reg, col_reg}<22'b0111110110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110110101000000010) && ({row_reg, col_reg}<22'b0111110110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110110101010000010) && ({row_reg, col_reg}<22'b0111110110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110110110000101101) && ({row_reg, col_reg}<22'b0111110111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110111000001010111) && ({row_reg, col_reg}<22'b0111110111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110111001000000010) && ({row_reg, col_reg}<22'b0111110111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110111001010000010) && ({row_reg, col_reg}<22'b0111110111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110111010000101101) && ({row_reg, col_reg}<22'b0111110111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111110111100001010111) && ({row_reg, col_reg}<22'b0111110111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111110111101000000010) && ({row_reg, col_reg}<22'b0111110111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111110111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111110111101010000010) && ({row_reg, col_reg}<22'b0111110111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111110111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111110111110000101101) && ({row_reg, col_reg}<22'b0111111000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111000000001010111) && ({row_reg, col_reg}<22'b0111111000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111000001000000010) && ({row_reg, col_reg}<22'b0111111000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111000001010000010) && ({row_reg, col_reg}<22'b0111111000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111000010000101101) && ({row_reg, col_reg}<22'b0111111000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111000100001010111) && ({row_reg, col_reg}<22'b0111111000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111000101000000010) && ({row_reg, col_reg}<22'b0111111000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111000101010000010) && ({row_reg, col_reg}<22'b0111111000110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111000110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111000110000101101) && ({row_reg, col_reg}<22'b0111111001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111001000001010111) && ({row_reg, col_reg}<22'b0111111001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111001001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111001001000000010) && ({row_reg, col_reg}<22'b0111111001001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111001001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111001001010000010) && ({row_reg, col_reg}<22'b0111111001010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111001010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111001010000101101) && ({row_reg, col_reg}<22'b0111111001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111001100001010111) && ({row_reg, col_reg}<22'b0111111001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111001101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111001101000000010) && ({row_reg, col_reg}<22'b0111111001101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111001101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111001101010000010) && ({row_reg, col_reg}<22'b0111111001110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111001110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111001110000101101) && ({row_reg, col_reg}<22'b0111111010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111010000001010111) && ({row_reg, col_reg}<22'b0111111010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111010001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111111010001000000010) && ({row_reg, col_reg}<22'b0111111010001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111010001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111010001010000010) && ({row_reg, col_reg}<22'b0111111010010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111010010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111010010000101101) && ({row_reg, col_reg}<22'b0111111010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111010100001010111) && ({row_reg, col_reg}<22'b0111111010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111010101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111111010101000000010) && ({row_reg, col_reg}<22'b0111111010101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111010101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111010101010000010) && ({row_reg, col_reg}<22'b0111111010110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111010110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111010110000101101) && ({row_reg, col_reg}<22'b0111111011000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111011000001010111) && ({row_reg, col_reg}<22'b0111111011001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111011001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111111011001000000010) && ({row_reg, col_reg}<22'b0111111011001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111011001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111011001010000010) && ({row_reg, col_reg}<22'b0111111011010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111011010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111011010000101101) && ({row_reg, col_reg}<22'b0111111011100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111011100001010111) && ({row_reg, col_reg}<22'b0111111011101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111011101000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111111011101000000010) && ({row_reg, col_reg}<22'b0111111011101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111011101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111011101010000010) && ({row_reg, col_reg}<22'b0111111011110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111011110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111011110000101101) && ({row_reg, col_reg}<22'b0111111100000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111100000001010111) && ({row_reg, col_reg}<22'b0111111100001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111100001000000001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=22'b0111111100001000000010) && ({row_reg, col_reg}<22'b0111111100001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111100001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111100001010000010) && ({row_reg, col_reg}<22'b0111111100010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111100010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111100010000101101) && ({row_reg, col_reg}<22'b0111111100100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111100100001010111) && ({row_reg, col_reg}<22'b0111111100101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111100101000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111111100101000000010) && ({row_reg, col_reg}<22'b0111111100101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111100101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111100101010000010) && ({row_reg, col_reg}<22'b0111111100110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111100110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111100110000101101) && ({row_reg, col_reg}<22'b0111111101000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111101000001010111) && ({row_reg, col_reg}<22'b0111111101001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111101001000000001)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b0111111101001000000010) && ({row_reg, col_reg}<22'b0111111101001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111101001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111101001010000010) && ({row_reg, col_reg}<22'b0111111101010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111101010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111101010000101101) && ({row_reg, col_reg}<22'b0111111101100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111101100001010111) && ({row_reg, col_reg}<22'b0111111101101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111101101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111101101000000010) && ({row_reg, col_reg}<22'b0111111101101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111101101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111101101010000010) && ({row_reg, col_reg}<22'b0111111101110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111101110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111101110000101101) && ({row_reg, col_reg}<22'b0111111110000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111110000001010111) && ({row_reg, col_reg}<22'b0111111110001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111110001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111110001000000010) && ({row_reg, col_reg}<22'b0111111110001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111110001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111110001010000010) && ({row_reg, col_reg}<22'b0111111110010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111110010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111110010000101101) && ({row_reg, col_reg}<22'b0111111110100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111110100001010111) && ({row_reg, col_reg}<22'b0111111110101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111110101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111110101000000010) && ({row_reg, col_reg}<22'b0111111110101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111110101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111110101010000010) && ({row_reg, col_reg}<22'b0111111110110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111110110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111110110000101101) && ({row_reg, col_reg}<22'b0111111111000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111111000001010111) && ({row_reg, col_reg}<22'b0111111111001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111111001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111111001000000010) && ({row_reg, col_reg}<22'b0111111111001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111111001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111111001010000010) && ({row_reg, col_reg}<22'b0111111111010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111111010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111111010000101101) && ({row_reg, col_reg}<22'b0111111111100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b0111111111100001010111) && ({row_reg, col_reg}<22'b0111111111101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111111101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b0111111111101000000010) && ({row_reg, col_reg}<22'b0111111111101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b0111111111101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b0111111111101010000010) && ({row_reg, col_reg}<22'b0111111111110000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b0111111111110000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b0111111111110000101101) && ({row_reg, col_reg}<22'b1000000000000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000000000001010111) && ({row_reg, col_reg}<22'b1000000000001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000000001000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000000000001000000010) && ({row_reg, col_reg}<22'b1000000000001010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000000001010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000000000001010000010) && ({row_reg, col_reg}<22'b1000000000010000101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000000010000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b1000000000010000101101) && ({row_reg, col_reg}<22'b1000000000100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000000100001010111) && ({row_reg, col_reg}<22'b1000000000101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000000101000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000000000101000000010) && ({row_reg, col_reg}<22'b1000000000101010000001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000000101010000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000000000101010000010) && ({row_reg, col_reg}<22'b1000000000110000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000000000110000101100) && ({row_reg, col_reg}<22'b1000000001000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000001000001010111) && ({row_reg, col_reg}<22'b1000000001001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000001001000000001)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=22'b1000000001001000000010) && ({row_reg, col_reg}<22'b1000000001001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000001001010000010) && ({row_reg, col_reg}<22'b1000000001010000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000000001010000101100) && ({row_reg, col_reg}<22'b1000000001100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000001100001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000000001100001011000) && ({row_reg, col_reg}<22'b1000000001101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000001101000000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b1000000001101000000010) && ({row_reg, col_reg}<22'b1000000001101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000001101010000010) && ({row_reg, col_reg}<22'b1000000001110000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000000001110000101100) && ({row_reg, col_reg}<22'b1000000010000001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000010000001010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000000010000001011000) && ({row_reg, col_reg}<22'b1000000010001000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000010001000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000000010001000000010) && ({row_reg, col_reg}<22'b1000000010001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000010001010000010) && ({row_reg, col_reg}<22'b1000000010010000101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000000010010000101100) && ({row_reg, col_reg}<22'b1000000010100001010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000010100001010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b1000000010100001011000) && ({row_reg, col_reg}<22'b1000000010101000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b1000000010101000000001) && ({row_reg, col_reg}<22'b1000000010101010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000010101010000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b1000000010101010000011) && ({row_reg, col_reg}<22'b1000000010110000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000010110000101011)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=22'b1000000010110000101100) && ({row_reg, col_reg}<22'b1000000011000001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000011000001011000) && ({row_reg, col_reg}<22'b1000000011001000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000011001000000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000000011001000000001) && ({row_reg, col_reg}<22'b1000000011001010000010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000011001010000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b1000000011001010000011) && ({row_reg, col_reg}<22'b1000000011010000101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000011010000101011)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=22'b1000000011010000101100) && ({row_reg, col_reg}<22'b1000000011100001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000011100001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000000011100001011001) && ({row_reg, col_reg}<22'b1000000011101000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000011101000000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b1000000011101000000001) && ({row_reg, col_reg}<22'b1000000011101010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000011101010000011) && ({row_reg, col_reg}<22'b1000000011110000101011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000000011110000101011) && ({row_reg, col_reg}<22'b1000000100000001011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000100000001011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b1000000100000001011001) && ({row_reg, col_reg}<22'b1000000100001000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b1000000100001000000000) && ({row_reg, col_reg}<22'b1000000100001010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000100001010000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000000100001010000100) && ({row_reg, col_reg}<22'b1000000100010000101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000100010000101010)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=22'b1000000100010000101011) && ({row_reg, col_reg}<22'b1000000100100001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000100100001011001) && ({row_reg, col_reg}<22'b1000000100100111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000100100111111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b1000000100101000000000) && ({row_reg, col_reg}<22'b1000000100101010000011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000100101010000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b1000000100101010000100) && ({row_reg, col_reg}<22'b1000000100110000101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000100110000101010)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=22'b1000000100110000101011) && ({row_reg, col_reg}<22'b1000000101000001011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000101000001011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000000101000001011010) && ({row_reg, col_reg}<22'b1000000101000111111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b1000000101000111111111) && ({row_reg, col_reg}<22'b1000000101001010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000101001010000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=22'b1000000101001010000101) && ({row_reg, col_reg}<22'b1000000101010000101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000101010000101001)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=22'b1000000101010000101010) && ({row_reg, col_reg}<22'b1000000101100001011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000101100001011010) && ({row_reg, col_reg}<22'b1000000101100111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000101100111111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b1000000101100111111111) && ({row_reg, col_reg}<22'b1000000101101010000100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000101101010000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000000101101010000101) && ({row_reg, col_reg}<22'b1000000101110000101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000101110000101001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b1000000101110000101010) && ({row_reg, col_reg}<22'b1000000110000001011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000110000001011010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b1000000110000001011011) && ({row_reg, col_reg}<22'b1000000110000111111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=22'b1000000110000111111110) && ({row_reg, col_reg}<22'b1000000110001010000101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000110001010000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b1000000110001010000110) && ({row_reg, col_reg}<22'b1000000110010000101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000110010000101000)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=22'b1000000110010000101001) && ({row_reg, col_reg}<22'b1000000110100001011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000110100001011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b1000000110100001011100) && ({row_reg, col_reg}<22'b1000000110100111111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000110100111111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000000110100111111110) && ({row_reg, col_reg}<22'b1000000110101010000110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000110101010000110) && ({row_reg, col_reg}<22'b1000000110110000101000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000000110110000101000) && ({row_reg, col_reg}<22'b1000000111000001011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000111000001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000000111000001011101) && ({row_reg, col_reg}<22'b1000000111000111111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000111000111111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b1000000111000111111101) && ({row_reg, col_reg}<22'b1000000111001010000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=22'b1000000111001010000111) && ({row_reg, col_reg}<22'b1000000111010000100111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000000111010000100111) && ({row_reg, col_reg}<22'b1000000111100001011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000111100001011101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b1000000111100001011110) && ({row_reg, col_reg}<22'b1000000111100111111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000111100111111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000000111100111111100) && ({row_reg, col_reg}<22'b1000000111101010000111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000000111101010000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000000111101010001000) && ({row_reg, col_reg}<22'b1000000111110000100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000000111110000100110)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=22'b1000000111110000100111) && ({row_reg, col_reg}<22'b1000001000000001011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001000000001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000001000000001011111) && ({row_reg, col_reg}<22'b1000001000000111111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001000000111111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000001000000111111011) && ({row_reg, col_reg}<22'b1000001000001010001000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001000001010001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000001000001010001001) && ({row_reg, col_reg}<22'b1000001000010000100101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=22'b1000001000010000100101) && ({row_reg, col_reg}<22'b1000001000100001011111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001000100001011111)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=22'b1000001000100001100000) && ({row_reg, col_reg}<22'b1000001000100111111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001000100111111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=22'b1000001000100111111010) && ({row_reg, col_reg}<22'b1000001000101010001010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001000101010001010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b1000001000101010001011) && ({row_reg, col_reg}<22'b1000001000110000100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001000110000100011)) color_data = 12'b011001100110;

		if(({row_reg, col_reg}>=22'b1000001000110000100100) && ({row_reg, col_reg}<22'b1000001001000001100000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001001000001100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b1000001001000001100001) && ({row_reg, col_reg}<22'b1000001001000111110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001001000111110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000001001000111111000) && ({row_reg, col_reg}<22'b1000001001001010001011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001001001010001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000001001001010001100) && ({row_reg, col_reg}<22'b1000001001010000100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001001010000100010)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b1000001001010000100011) && ({row_reg, col_reg}<22'b1000001001100001100010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001001100001100010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=22'b1000001001100001100011) && ({row_reg, col_reg}<22'b1000001001100111110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001001100111110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==22'b1000001001100111110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=22'b1000001001100111110111) && ({row_reg, col_reg}<22'b1000001001101010001101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001001101010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=22'b1000001001101010001110) && ({row_reg, col_reg}<22'b1000001001110000100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001001110000100000)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=22'b1000001001110000100001) && ({row_reg, col_reg}<22'b1000001010000001100100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001010000001100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b1000001010000001100101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=22'b1000001010000001100110) && ({row_reg, col_reg}<22'b1000001010000111110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001010000111110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b1000001010000111110100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000001010000111110101) && ({row_reg, col_reg}<22'b1000001010001010001111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001010001010001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=22'b1000001010001010010000) && ({row_reg, col_reg}<22'b1000001010010000011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001010010000011110)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=22'b1000001010010000011111) && ({row_reg, col_reg}<22'b1000001010100001100111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001010100001100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==22'b1000001010100001101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==22'b1000001010100001101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000001010100001101010) && ({row_reg, col_reg}<22'b1000001010100111101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001010100111101110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==22'b1000001010100111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b1000001010100111110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b1000001010100111110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=22'b1000001010100111110010) && ({row_reg, col_reg}<22'b1000001010101010010010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==22'b1000001010101010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==22'b1000001010101010010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b1000001010101010010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=22'b1000001010101010010101) && ({row_reg, col_reg}<22'b1000001010110000011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==22'b1000001010110000011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==22'b1000001010110000011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==22'b1000001010110000011011)) color_data = 12'b101010101010;





































































		if(({row_reg, col_reg}>=22'b1000001010110000011100) && ({row_reg, col_reg}<=22'b1000101100110001110101)) color_data = 12'b000000001111;
	end
endmodule